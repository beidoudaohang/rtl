//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : pixelformat_sel
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/12/5 14:17:37	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ͼ��ѡ��ģ��
//              1)  : MT9P031ʱ����ģ��û�������ã�Ϊ���Ժ����չ����ƣ�������ģ��
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module pixelformat_sel # (
	parameter				SENSOR_DAT_WIDTH	= 10	,	//sensor ���ݿ��
	parameter				REG_WD				= 32		//�Ĵ���λ��
	)
	(
	//Sensor�����ź�
	input								clk				,	//����ʱ��
	input								i_fval			,	//���ź�
	input								i_lval			,	//���ź�
	input	[SENSOR_DAT_WIDTH-1:0]		iv_pix_data		,	//ͼ������
	//�Ĵ�������
	input	[REG_WD-1:0]				iv_pixel_format	,	//0x01080001:Mono8��0x01100003:Mono10��0x01080008:BayerGR8��0x0110000C:BayerGR10
	//ͼ�����
	output								o_fval			,	//����Ч
	output								o_lval			,	//����Ч
	output	[SENSOR_DAT_WIDTH-1:0]		ov_pix_data			//ͼ������
	);

	//	ref signals



	//	ref ARCHITECTURE

	assign	o_fval		= i_fval;
	assign	o_lval		= i_lval;
	assign	ov_pix_data	= iv_pix_data;


endmodule