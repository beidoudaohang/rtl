//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : dcm_pix
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/2/28 13:11:28	:|  ��ʼ�汾
//  -- ��  ǿ       :| 2015/12/21 14:40:20	:|  mer_230_060u3x���36MHzʱ��
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module dcm_pix (
	input         clk_in		,	//ʱ������
	input         dcm_reset		,	//DCM��λ������Ч
	output        clk_fx_out	,	//clkfx���
	output        clk_fxdv_out	,	//clkfx���
	output        locked			//DCM����������Ч
	);

	//	ref signals
	wire 				clkfx			;
	wire 				clkfxdv			;

	//	ref ARCHITECTURE

	//  -------------------------------------------------------------------------------------
	//	dcm ����
	//  -------------------------------------------------------------------------------------
	DCM_CLKGEN # (
	.CLKFXDV_DIVIDE        (2				),
	.CLKFX_DIVIDE          (4				),
	.CLKFX_MULTIPLY        (11				),
	.SPREAD_SPECTRUM       ("NONE"			),
	.STARTUP_WAIT          ("FALSE"			),
	.CLKIN_PERIOD          (25.000			),
	.CLKFX_MD_MAX          (0.000			)
	)
	DCM_CLKGEN_inst (
	// Input clock
	.CLKIN                 (clk_in			),
	// Output clocks
	.CLKFX                 (clkfx			),
	.CLKFX180              (				),
	.CLKFXDV               (clkfxdv			),
	// Ports for dynamic reconfiguration
	.PROGCLK               (1'b0			),
	.PROGDATA              (1'b0			),
	.PROGEN                (1'b0			),
	.PROGDONE              (				),
	// Other control and status signals
	.FREEZEDCM             (1'b0			),
	.LOCKED                (locked			),
	.STATUS                (				),
	.RST                   (dcm_reset		)
	);

	//  -------------------------------------------------------------------------------------
	//	clkfxȫ������
	//  -------------------------------------------------------------------------------------
	BUFGCE clkfx_buf (
	.I						(clkfx			),
	.CE						(locked			),
	.O						(clk_fx_out		)
	);

	//  -------------------------------------------------------------------------------------
	//	clkfxdvȫ������
	//  -------------------------------------------------------------------------------------
	BUFGCE clkfxdv_buf (
	.I						(clkfxdv		),
	.CE						(locked			),
	.O						(clk_fxdv_out	)
	);


endmodule
