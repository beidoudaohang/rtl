//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : testcase_1
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/4/10 16:50:28	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ���ڴ�С��16x16�������ź���Ч������ģʽ�µ�����״��
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module testcase_1 ();

	//	ref signals
	//	===============================================================================================
	//	--ref parameter
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	TESTCASE
	//	-------------------------------------------------------------------------------------
	parameter	TESTCASE_NUM			= "testcase_1"			;	//����ģ����Ҫʹ���ַ���
	//	-------------------------------------------------------------------------------------
	//	sensor model parameter
	//	-------------------------------------------------------------------------------------
	parameter	PYTHON_IMAGE_SRC				= "RANDOM"			;	//"RANDOM" or "FILE" or "LINE_INC" or "FRAME_INC" or "FRAME_INC_NO_RST" or "PIX_INC_NO_FVAL" or "PIX_INC"
	parameter	PYTHON_DATA_WIDTH				= 10				;	//���ݿ��
	parameter	PYTHON_SOURCE_FILE_PATH			= "source_file/"	;	//����Դ�ļ�·��
	parameter	PYTHON_GEN_FILE_EN				= 0					;	//0-���ɵ�ͼ��д���ļ���1-���ɵ�ͼ��д���ļ�
	parameter	PYTHON_GEN_FILE_PATH			= "gen_file/"		;	//����������Ҫд���·��
	parameter	PYTHON_NOISE_EN					= 0					;	//0-������������1-��������

	//	-------------------------------------------------------------------------------------
	//	dut paramter
	//	-------------------------------------------------------------------------------------
	parameter	SER_FIRST_BIT		= "MSB"	;
	parameter	END_STYLE			= "LITTLE"	;
	parameter	SER_DATA_RATE		= "DDR"	;
	parameter	DESER_CLOCK_ARC		= "BUFPLL"	;
	parameter	CHANNEL_NUM			= 4	;
	parameter	DESER_WIDTH			= 5	;
	parameter	CLKIN_PERIOD_PS		= 3030	;
	parameter	DATA_DELAY_TYPE		= "DIFF_PHASE_DETECTOR"	;
	parameter	DATA_DELAY_VALUE	= 0	;
	parameter	BITSLIP_ENABLE		= "TRUE"	;

	//	-------------------------------------------------------------------------------------
	//	monitor paramter
	//	-------------------------------------------------------------------------------------


	//	-------------------------------------------------------------------------------------
	//	testcase parameter
	//	-------------------------------------------------------------------------------------
	parameter	CLK_PERIOD				= 20	;	//ʱ��Ƶ�ʣ�50MHz

	//	===============================================================================================
	//	--ref signal
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	sensor signal
	//	-------------------------------------------------------------------------------------
	reg					clk_python		= 1'b0;

	//	-------------------------------------------------------------------------------------
	//	dut signal
	//	-------------------------------------------------------------------------------------
	wire								i_clk_p	;
	wire								i_clk_n	;
	wire	[CHANNEL_NUM:0]				iv_data_p	;
	wire	[CHANNEL_NUM:0]				iv_data_n	;
	wire								reset	;
	reg									i_bitslip_en	;

	//	ref ARCHITECTURE

	//	===============================================================================================
	//	ref ***tb ��ģ�鼤��***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	--ref Sensor
	//	-------------------------------------------------------------------------------------
	always	#(CLK_PERIOD/2.0)	clk_python	= !clk_python;



	//	-------------------------------------------------------------------------------------
	//	--ref DUT
	//	-------------------------------------------------------------------------------------
	assign	i_clk_p					= driver_python.o_clk_p;
	assign	i_clk_n					= driver_python.o_clk_n;
	assign	iv_data_p				= {driver_python.ov_data_p,driver_python.o_ctrl_p};
	assign	iv_data_n				= {driver_python.ov_data_n,driver_python.o_ctrl_n};

	assign	reset					= 1'b0;

	//	-------------------------------------------------------------------------------------
	//	--ref ����ʱ��
	//	-------------------------------------------------------------------------------------
	initial begin
		#200
		#20000
		$stop;
	end

	initial begin
		//$display("** ");
		//#1000000
		i_bitslip_en	= 1'b1;
		#2520
		i_bitslip_en	= 1'b0;
	end


	//	===============================================================================================
	//	ref ***����bfm task***
	//	===============================================================================================



endmodule
