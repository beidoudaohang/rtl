//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : data_align
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/12/5 15:44:31	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ����ƴ��ģ��
//              1)  : ����pixel format������λ��ѡ��ƴ�ӷ�ʽ�����λ��̶�Ϊ32bit
//
//              2)  : ���pixel format������λ����8bit��ѡ���������ݵĸ�8bit��ÿ4������ƴ��Ϊ1��32bit���ݣ��ȵ��������ݷ��ڵ�λ
//
//              3)  : ���pixel format������λ����10bit��ѡ���������ݸ�10bit��ÿ2������ƴ��Ϊ1��32bit���ݣ��ȵ��������ݷ��ڵ�λ
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module data_align # (
	parameter	SENSOR_DAT_WIDTH	= 10	,	//sensor ���ݿ��
	parameter	REG_WD				= 32	,	//�Ĵ���λ��
	parameter	DATA_WD				= 32		//�����������λ������ʹ��ͬһ���
	)
	(
	//Sensor�����ź�
	input								clk				,	//����ʱ��
	input								i_fval			,	//���ź�
	input								i_lval			,	//���ź�
	input	[SENSOR_DAT_WIDTH-1:0]		iv_pix_data		,	//ͼ������
	//�Ҷ�ͳ����ؼĴ���
	input	[REG_WD-1:0]				iv_pixel_format	,	//���ظ�ʽ�Ĵ�����0x01080001:Mono8��0x01100003:Mono10��0x01080008:BayerGR8��0x0110000C:BayerGR10
	//���
	output								o_fval			,	//����Ч
	output								o_pix_data_en	,	//������Ч�źţ�����ƴ��֮���ʹ���źţ��൱��ʱ�ӵ�2��Ƶ����4��Ƶ
	output	[DATA_WD-1:0]				ov_pix_data			//ͼ������
	);

	//	ref signals
	reg							format8_sel		= 1'b0;
	reg		[DATA_WD-1:0]		pix_data_shift	= {DATA_WD{1'b0}};
	reg		[DATA_WD-1:0]		pix_data_reg	= {DATA_WD{1'b0}};
	reg		[1:0]				pix_cnt			= 2'b0;
	reg							data_en			= 1'b0;
	reg							data_en_dly		= 1'b0;
	reg							fval_dly0		= 1'b0;
	reg							fval_dly1		= 1'b0;

	//	ref ARCHITECTURE
	//  ===============================================================================================
	//	ref ***�ж����ݸ�ʽ***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	Mono8		- 0x01080001	-> 0x1081	-> 0001,0000,1000,,,,0001
	//	Mono10		- 0x01100003	-> 0x1103	-> 0001,0001,0000,,,,0011
	//	BayerGR8	- 0x01080008	-> 0x1088	-> 0001,0000,1000,,,,1000
	//	BayerGR10	- 0x0110000C	-> 0x110C	-> 0001,0001,0000,,,,1100
	//											   --------!-!-------!!!!
	//                                                     ^    ^       ^------bit0
	//                                             bit20---|    |---bit16
	//	����� ! �ģ����ǲ���Ƚϵ�bit.�ֱ��� bit 20 19 3-0
	//  -------------------------------------------------------------------------------------
	//  -------------------------------------------------------------------------------------
	//	format8_sel
	//	1.�ж����ظ�ʽ�Ƿ�ѡ��8bit���ظ�ʽ
	//	2.ʹ��6bit�ж�����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		case({iv_pixel_format[20],iv_pixel_format[19],iv_pixel_format[3:0]})
			6'b010001	: format8_sel	<= 1'b1;
			6'b011000	: format8_sel	<= 1'b1;
			default		: format8_sel	<= 1'b0;
		endcase
	end

	//  ===============================================================================================
	//	ref ***������λ***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	������λ�Ĵ���
	//	1.��������ʱ����λ�Ĵ�������
	//	2.������Ч������Чʱ��������ظ�ʽ��8bit��ÿ������ռ��1��byte��ֻȡ���صĸ�8bit
	//	3.������Ч������Чʱ��������ظ�ʽ��10bit��ÿ������ռ��2��byte����ֻȡ���صĸ�10bit����λ���0
	//	4.������λ�Ĵ���λ��-32bit
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!i_fval) begin
			pix_data_shift	<= {DATA_WD{1'b0}};
		end
		else begin
			if(i_lval) begin
				//  -------------------------------------------------------------------------------------
				//	���ظ�ʽ8bit
				//  -------------------------------------------------------------------------------------
				if(format8_sel) begin
					pix_data_shift	<= {iv_pix_data[SENSOR_DAT_WIDTH-1:SENSOR_DAT_WIDTH-8],pix_data_shift[DATA_WD-1:8]};
				end
				//  -------------------------------------------------------------------------------------
				//	���ظ�ʽ10bit
				//  -------------------------------------------------------------------------------------
				else begin
					pix_data_shift	<= {6'b0,iv_pix_data[SENSOR_DAT_WIDTH-1:SENSOR_DAT_WIDTH-10],pix_data_shift[DATA_WD-1:16]};
				end
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	���ؼ�����
	//	1.������ʱ������
	//	2.����Ч������Чʱ���������ۼ�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!i_fval) begin
			pix_cnt	<= 2'b0;
		end
		else begin
			if(i_lval) begin
				pix_cnt	<= pix_cnt + 1'b1;
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	data_en ����ʹ���źţ�����o_lval
	//	1.����������ʱ������ʹ�ܱ�����0.
	//	2.������Ч��ʱ�򣬵�����Чʱ��������ظ�ʽ8bit��ÿ4�����ڣ�����1������ʹ��
	//	3.������Ч��ʱ�򣬵�����Чʱ��������ظ�ʽ10bit��ÿ2�����ڣ�����1������ʹ��
	//	4.������Ч��ʱ�򣬵�����Чʱ������ʹ����Ч
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!i_fval) begin
			data_en	<= 1'b0;
		end
		else begin
			if(i_lval) begin
				//  -------------------------------------------------------------------------------------
				//	���ظ�ʽ8bit
				//  -------------------------------------------------------------------------------------
				if(format8_sel) begin
					if(pix_cnt==2'b11) begin
						data_en	<= 1'b1;
					end
					else begin
						data_en	<= 1'b0;
					end
				end
				//  -------------------------------------------------------------------------------------
				//	���ظ�ʽ10bit
				//  -------------------------------------------------------------------------------------
				else begin
					if(pix_cnt[0]==1'b1) begin
						data_en	<= 1'b1;
					end
					else begin
						data_en	<= 1'b0;
					end
				end
			end
			else begin
				data_en	<= 1'b0;
			end
		end
	end

	//  ===============================================================================================
	//	ref ***�г��źš��������***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	fval ���
	//	1.�ӽ�β������������ʱ��2��ʱ����������Ҫ��fval��ʱ2��ʱ������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_dly0	<= i_fval;
		fval_dly1	<= fval_dly0;
	end

	//	-------------------------------------------------------------------------------------
	//	��data_en��ʱ1�ģ���Ϊ���ݵĴ����ͺ���һ�ģ�����Ҫ��ʱ
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		data_en_dly	<= data_en;
	end

	//	-------------------------------------------------------------------------------------
	//	�ж�������ݣ������ʹ�ܣ������Ϊȫ��
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(data_en) begin
			pix_data_reg	<= pix_data_shift;
		end
		else begin
			pix_data_reg	<= {DATA_WD{1'b0}};
		end
	end

	//  -------------------------------------------------------------------------------------
	//	���
	//  -------------------------------------------------------------------------------------
	assign	o_pix_data_en	= data_en_dly;
	assign	ov_pix_data		= pix_data_reg;
	assign	o_fval			= fval_dly1;



endmodule
