//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : dna
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/12/12 16:10:44	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ģ�����ʱ����clk_osc_bufg 40MHz��DNAģ�����ֻ��֧�ֵ�2MHz��Ƶ�ʣ������dnaģ���ڲ�
//					��clk_osc_bufg��ƵΪ1MHz��ʱ��-clk_dna����clk_dna����FPGA�ڲ���dnaģ�顣
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module dna # (
	parameter		LONG_REG_WD				= 64	,	//���Ĵ���λ��
	parameter		REG_INIT_VALUE			= "TRUE"	//�Ĵ����Ƿ��г�ʼֵ
	)
	(
	input						clk					,	//40MHz
	input						reset				,	//40MHz��λ�ź�
	output	[LONG_REG_WD-1:0]	ov_dna_reg			,	//clk_dnaʱ���򣬶���dna֮���ȶ�����
	input	[LONG_REG_WD-1:0]	iv_encrypt_reg		,	//clk_osc_bufgʱ����
	output						o_encrypt_state			//clk_dnaʱ���򣬼���״̬��1-���ܳɹ���0-����ʧ��
	);

	//	ref signals
	reg		[4:0]		clk_div_cnt		= 5'b0;
	wire				clk_dna			;
	reg		[6:0]		flow_cnt		= 7'b0;
	reg					dna_read		= 1'b0;
	reg					dna_shift		= 1'b0;
	reg		[56:0]		dna_reg			= 57'b0;
	reg		[55:0]		dna_enc_reg0	= 56'b0;
	wire	[63:0]		dna_enc_reg1	;
	reg					encrypt_state_reg	= 1'b0;


	//	ref ARCHITECTURE

	//  ===============================================================================================
	//	ref ***���� DNA ģ��***
	//	1.bit56�̶���1��bit55�̶���0��������ģ������ֻ��bit56�̶�Ϊ0��
	//	2.��read=1ʱ�����ڲ�����ת�Ƶ���λ�Ĵ����ϣ�ͬʱdout=bit56=1����shift=1ʱ����bit55�Ƶ�dout�ϡ����Ҫ��λ��57bit���ݣ�shiftֻ��56��ʱ�ӡ�
	//	3.ug380�涨����������£�SHIFT��clk=0������clk�½��أ���0��Ϊ1
	//  ===============================================================================================
	DNA_PORT # (
	.SIM_DNA_VALUE	(57'h043210000001234	)  // Specifies the Pre-programmed factory ID value
	)
	DNA_PORT_inst (
	.DOUT		(dna_dout	),	// 1-bit output: DNA output data
	.CLK		(clk_dna	),	// 1-bit input: Clock input
	.DIN		(1'b0		),	// 1-bit input: User data input pin
	.READ		(dna_read	),	// 1-bit input: Active high load DNA, active low read input
	.SHIFT		(dna_shift	)	// 1-bit input: Active high shift enable input
	);

	//  ===============================================================================================
	//	ref ***��DNA_PORT���߼�***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	��Ƶ������
	//	1.40MHz 32 ��Ƶ��1.25MHz
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(reset) begin
			clk_div_cnt	<= 5'b0;
		end
		else begin
			clk_div_cnt	<= clk_div_cnt + 1'b1;
		end
	end
	assign	clk_dna	= clk_div_cnt[4];

	//  -------------------------------------------------------------------------------------
	//	�� dna ���̿��Ƶļ�����
	//	1.��clk dna�½��ص�ʱ��flow cnt����
	//	2.��flow cnt bit6=1 �����ӵ�64ʱ��ֹͣ
	//  ------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(reset) begin
			flow_cnt	<= 7'b0;
		end
		else begin
			//��ʱclk dna�����½���
			if(clk_div_cnt==5'h1f) begin
				if(flow_cnt[6]) begin
					flow_cnt	<= flow_cnt;
				end
				else begin
					flow_cnt	<= flow_cnt + 1'b1;
				end
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	�������źţ�ʹ dna_port �е�����ת�Ƶ���λ�Ĵ�������
	//	1.read�ź���clk dna���½��ض��룬�ο�ug382��shift��Լ��
	//  ------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(flow_cnt==7'd2) begin
			dna_read	<= 1'b1;
		end
		else begin
			dna_read	<= 1'b0;
		end
	end

	//  -------------------------------------------------------------------------------------
	//	������λ�ź�
	//	1.shift�ź���clk dna���½��ض��룬Ϊ���Ƿ���ug380�Ĺ涨
	//	2.shift�źſ����56��ʱ������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(flow_cnt>=7'd3 && flow_cnt<=7'd58) begin
			dna_shift	<= 1'b1;
		end
		else begin
			dna_shift	<= 1'b0;
		end
	end

	//  -------------------------------------------------------------------------------------
	//	���� dna ģ�����������
	//	1.��read=1ʱ��dou���1����dna_data�����bit
	//	2.��read=0 shift=1ʱ����ʼ��λ
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(flow_cnt>=7'd2 && flow_cnt<=7'd58) begin
			//��ʱclk dna�����½���
			if(clk_div_cnt==5'h1f) begin
				dna_reg	<= {dna_reg[55:0],dna_dout};
			end
		end
	end
	assign	ov_dna_reg	= {7'b0,dna_reg};

	//  ===============================================================================================
	//	ref ***�����㷨***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	���ɼ�����
	//	1.��dna����֮�󣬵�7���ֽڰ�λ����0xaa
	//	2.����ֽ���0x47����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(flow_cnt[6]) begin
			dna_enc_reg0	<= dna_reg[55:0] & 56'haaaaaa_aaaaaaaa;
		end
		else begin
			dna_enc_reg0	<= 56'h0;
		end
	end
	assign	dna_enc_reg1	= {8'h47,dna_enc_reg0};

	//  -------------------------------------------------------------------------------------
	//	�жϼ���״̬
	//	1.����̼����õļ�������fpga�����ļ�����һ���������ͨ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(dna_enc_reg1==iv_encrypt_reg) begin
			encrypt_state_reg	<= 1'b1;
		end
		else begin
			encrypt_state_reg	<= 1'b0;
		end
	end

	generate
		if(REG_INIT_VALUE=="TRUE") begin
			assign	o_encrypt_state	= 1'b1;
		end
		else begin
			assign	o_encrypt_state	= encrypt_state_reg;
		end
	endgenerate





endmodule