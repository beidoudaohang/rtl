//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : mer_1810_21u3x
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����     :|  �޸�˵��
//---------------------------------------------------------------------------------------
//  -- ��ǿ         :| 2014/11/25   :|  ���������ź�����
//	-- �Ϻ���		:| 2015/3/30 	:|	��д��Ķ���ģ�����Ͻ���
//	-- �Ϻ���		:| 2015/9/23  	:|	��mer-500-14u3x��ֲ��mer-1520-13u3x
//	-- �ܽ�		:| 2016/3/23   	:|	��mer-1520-13u3x��ֲ��mer-1820-20u3x
//	-- �Ϻ���		:| 2016/6/23   	:|	�������ָ��� ��Ϊ mer-1810-21u3x
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1) 	: ��ģ����mer����1820����20u3x����Ķ���ģ�飬��Ҫ������xxxx����ģ��
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------
module mer_1810_21u3x  # (
	//  ===============================================================================================
	//	ref �ⲿ��������
	//	----��Ϊ parameter �Ĳ��������ⲿ�ӿ���أ�����ⲿ�ӿ��иĶ�����ô���������Ӧ����
	//  ===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	Sensor��ز���
	//	-------------------------------------------------------------------------------------
	parameter	SENSOR_DAT_WIDTH			= 12					,	//Sensor ���ݿ��
	parameter	PHY_NUM						= 2						,	//HiSPi PHY������
	parameter	PHY_CH_NUM					= 4						,	//ÿ·HiSPi PHY������ͨ����
	parameter	PIX_CLK_FREQ_KHZ			= 55000					,	//����ʱ��Ƶ�ʣ���λKHZ���ܶ�ģ���ø�ʱ����Ϊ��ʱ������˱���д������ʱ�ӵ�Ƶ��
	parameter	BAYER_PATTERN				= "GR"					,	//"GR" "RG" "GB" "BG"
	parameter	SENSOR_MAX_WIDTH			= 4912					,	//Sensor��������Ч��ȣ�������ʱ��Ϊ��λ
	parameter	SENSOR_MAX_HEIGHT			= 3684					,	//Sensor������Ч�и���������Ϊ��λ
	parameter	SHORT_LINE_LENGTH_PCK		= 5568					,	//sensor������������ֵ�����ֵ��д��sensor�Ĵ�����ʮ���Ʊ�ʾ
	//	-------------------------------------------------------------------------------------
	//	�⴮��صĲ���
	//	-------------------------------------------------------------------------------------
	parameter	DIFF_TERM					= "TRUE"				,	//Differential Termination
	parameter	IOSTANDARD					= "LVDS_33"				,	//Specifies the I/O standard for this buffer
	parameter	SER_FIRST_BIT				= "LSB"					,	//"LSB" or "MSB" , first bit to the receiver
	parameter	END_STYLE					= "LITTLE"				,	//"LITTLE" or "BIG" , "LITTLE" - {CHANNEL3 CHANNE2 CHANNEL1 CHANNEL0}. "BIG" - {CHANNEL0 CHANNEL1 CHANNEL2 CHANNEL3}.
	parameter	SER_DATA_RATE				= "DDR"					,	//"DDR" or "SDR" ����Ĵ���ʱ�Ӳ�����ʽ
	parameter	DESER_CLOCK_ARC				= "BUFPLL"				,	//"BUFPLL" or "BUFIO2" , deserializer clock achitecture
	parameter	DESER_WIDTH					= 6						,	//ÿ��ͨ���⴮��� 2-8
	parameter	CLKIN_PERIOD_PS				= 3030					,	//����ʱ��Ƶ�ʣ�PSΪ��λ��ֻ��BUFPLL��ʽ�����á�
	parameter	DATA_DELAY_TYPE				= "DIFF_PHASE_DETECTOR"	,	//"DEFAULT", "DIFF_PHASE_DETECTOR", "FIXED", "VARIABLE_FROM_HALF_MAX", "VARIABLE_FROM_ZERO"
	parameter	DATA_DELAY_VALUE			= 0						,	//0-255������ܳ��� 1 UI
	parameter	BITSLIP_ENABLE				= "FALSE"				,	//"TRUE" "FALSE" iserdes �ֱ߽���빦��
	parameter	PLL_RESET_SIMULATION		= "FALSE"				,	//�⴮PLL��λ��ʹ�ܷ���ģʽ����λʱ���̣����ٷ���
	//	-------------------------------------------------------------------------------------
	//	DDR3�Ĳ���
	//	-------------------------------------------------------------------------------------
	parameter	NUM_DQ_PINS					= 16 				,	//DDR3���ݿ��
	parameter	MEM_ADDR_WIDTH				= 13 				,	//DDR3��ַ���
	parameter	MEM_BANKADDR_WIDTH			= 3  				,	//DDR3bank���
	parameter	DDR3_MEMCLK_FREQ			= 320				,	//DDR3ʱ��Ƶ��
	parameter	MEM_ADDR_ORDER				= "ROW_BANK_COLUMN"	,	//DDR3��ַ�Ų�˳��
	parameter 	DDR3_RST_ACT_LOW          	= 0					,   // # = 1 for active low reset,# = 0 for active high reset.
	parameter	DDR3_MEM_DENSITY			= "1Gb"				,	//DDR3����
	parameter	DDR3_TCK_SPEED				= "15E"				,	//DDR3���ٶȵȼ�
	parameter	DDR3_SIMULATION				= "FALSE"			,	//�򿪷�����Լ��ٷ����ٶȣ�����ʵ�ʲ��ֲ���ʱ�����ܴ򿪷��档
	parameter	DDR3_P0_MASK_SIZE			= 8					,	//p0��mask size
	parameter	DDR3_P1_MASK_SIZE			= 8					,	//p1��mask size
	parameter	DDR3_CALIB_SOFT_IP			= "TRUE"			,	//����ʱ�����Բ�ʹ��У׼�߼�
	//	-------------------------------------------------------------------------------------
	//	GPIF����λ��
	//	-------------------------------------------------------------------------------------
	parameter	GPIF_DAT_WIDTH				= 32				,	//GPIF���ݿ��
	//	-------------------------------------------------------------------------------------
	//	GPIO��������λ�����ڴ���
	//	-------------------------------------------------------------------------------------
	parameter	NUM_GPIO					= 2						//GPIO����
	)
	(
	//  ===============================================================================================
	//  ��һ���֣�����ʱ���ź�
	//  ===============================================================================================
	input									clk_osc				,	//�������ţ�40MHz�����ⲿ����
	//  ===============================================================================================
	//  �ڶ����֣�sensor�ӿ��ź�
	//  ===============================================================================================
	input		[PHY_NUM-1:0]				pix_clk_p			,	//�������ţ�Sensor������330MHz��HiSpi���ʱ��
	input		[PHY_NUM-1:0]				pix_clk_n			,	//�������ţ�Sensor������330MHz��HiSpi���ʱ��
	input		[PHY_CH_NUM*PHY_NUM-1:0]	iv_pix_data_p		,	//�������ţ�Sensor������HiSPi������ݽӿ�
	input		[PHY_CH_NUM*PHY_NUM-1:0]	iv_pix_data_n		,	//�������ţ�Sensor������HiSPi������ݽӿ�
	input									i_sensor_strobe		,	//�������ţ�Sensor����������Ч��������ź�
	output									o_trigger			,	//������ţ�FPGA�����sensor�Ĵ����źţ�����Ч
	output									o_sensor_reset_n	,	//������ţ����ӵ�Sensor��Sensor�ĸ�λ�źţ�����Ч������1ms��FPGA������ɺ������������������в���λSensor
	output									o_clk_sensor		,	//Sensor��ʱ�ӣ�20Mhz����40M����������
	//  ===============================================================================================
	//  �ڶ����֣�GPIF�ӿ��ź�
	//  ===============================================================================================
	output									o_clk_usb_pclk		,	//������ţ����ӵ�3014��GPIF�ӿڵ�ʱ��100MHz��ʹ��ODDR�������FPGA �����ϣ�ʱ���½�����gpif���ݶ���
	output		[GPIF_DAT_WIDTH-1:0]		ov_usb_data			,	//������ţ����ӵ�3014��GPIF�ӿڵ����ݣ�clk_gpif ʱ������FPGA�����ϣ�o_clk_usb_pclk��ov_usb_data����
	output		[1:0]						ov_usb_fifoaddr		,	//������ţ����ӵ�3014��GPIF fifo��ַ��clk_gpif ʱ����00��11���棬��FPGA�����ϣ�o_clk_usb_pclk��ov_usb_data����
	output									o_usb_slwr_n		,	//������ţ����ӵ�3014��GPIF д�źţ�clk_gpif ʱ����
	output									o_usb_pktend_n		,	//������ţ����ӵ�3014��GPIF �������źţ�clk_gpif ʱ����
	input									i_usb_flagb_n		,	//�������ţ����ӵ�3014��3014������o_clk_usb_pclk ʱ����GPIF��ǰDMAbuffer���źţ��� clk_gpif ����λ���Ϊ���첽�źţ���Ҫ�� u3_interface ģ��������ʱ������
	//  ===============================================================================================
	//  �������֣�SPI�ӿ��ź�
	//  ===============================================================================================
	input									i_usb_spi_sck		,	//�������ţ�3014������SPIʱ�ӣ���������10Mhz���û�����463KhzƵ�ʣ�FPGA�趼���㡣���̼����û�����ʱ���ź�ռ�ձȿ��ܻ��нϴ�仯�����ź���С��ȱ�֤>384ns
	input									i_usb_spi_mosi		,	//�������ţ�3014������SPI�������룬�źſ�ȿ��ܻ��нϴ�仯�����ź���С��ȱ�֤>384ns
	input									i_spi_cs_n_fpga		,	//�������ţ�3014������SPI FPGAƬѡ���̼���һ���ܱ�ֻ֤�з���FPGAʱƬѡ�����ͣ�FPGA��Ҫ�����쳣��Ƭѡ
	output									o_usb_spi_miso		,	//������ţ����ӵ�3014���ⲿ��flash�����������SPI���������ֻ�ж�����ͨ��֮��������Ч���ݣ�������衣Ƭѡ��Чʱ����������
	//  ===============================================================================================
	//  ���Ĳ��֣�IO�ӿ��ź�
	//  ===============================================================================================
	input									i_optocoupler		,	//�������ţ�������������ȴ�0��������п��ܣ���������ë�̣���ȴ���֡����ʱ��Ҫ�����½��ص��󴥷����첽�ź�
	input		[NUM_GPIO-1:0]				iv_gpio				,	//�������ţ�������������˫��IO������ˣ���ȴ�0��������п��ܣ��������ܸ��ţ��첽�źš�˫��IO����Ϊ����ʱ������Ϊ0
	output									o_optocoupler		,	//������ţ����ӵ�������������·����ʱ��������ʱ7~44us��������ʱ9~35us
	output		[NUM_GPIO-1:0]				ov_gpio				,	//������ţ����ӵ������ܣ�˫��IO������ˣ���ʱ<1us,˫��IO����Ϊ����ʱ������Ϊ0
	output									o_f_led_gre			,	//������ţ����ӵ�LED����ɫָʾ�ƣ��ߵ�ƽ����
	output									o_f_led_red			,	//������ţ����ӵ�LED����ɫָʾ�ƣ��ߵ�ƽ����
	//  ===============================================================================================
	//  ���岿�֣�DDR3�ӿ��ź�
	//  ������ʹ���ź�����ddr3оƬ�ⲿ�ӿ��źţ������źŶ���ο���׼��ddr3�ӿ�
	//  ===============================================================================================
	inout  		[NUM_DQ_PINS-1:0]			mcb1_dram_dq		,	//DDR3������ţ������ź�
	output 		[MEM_ADDR_WIDTH-1:0]		mcb1_dram_a			,	//DDR3������ţ���ַ�ź�
	output 		[MEM_BANKADDR_WIDTH-1:0]	mcb1_dram_ba		,	//DDR3������ţ�Bank��ַ�ź�
	output									mcb1_dram_ras_n		,	//DDR3������ţ��е�ַѡͨ
	output									mcb1_dram_cas_n		,	//DDR3������ţ��е�ַѡͨ
	output									mcb1_dram_we_n		,	//DDR3������ţ�д�ź�
	output									mcb1_dram_odt		,	//DDR3������ţ��迹ƥ���ź�
	output									mcb1_dram_reset_n	,	//DDR3������ţ���λ�ź�
	output									mcb1_dram_cke		,	//DDR3������ţ�ʱ��ʹ���ź�
	output									mcb1_dram_dm		,	//DDR3������ţ����ֽ����������ź�
	inout 									mcb1_dram_udqs		,	//DDR3������ţ����ֽڵ�ַѡͨ�ź���
	inout 									mcb1_dram_udqs_n	,	//DDR3������ţ����ֽڵ�ַѡͨ�źŸ�
	inout 									mcb1_rzq			,	//DDR3������ţ�����У׼
	output									mcb1_dram_udm		,	//DDR3������ţ����ֽ����������ź�
	inout 									mcb1_dram_dqs		,	//DDR3������ţ����ֽ�����ѡͨ�ź���
	inout 									mcb1_dram_dqs_n		,	//DDR3������ţ����ֽ�����ѡͨ�źŸ�
	output									mcb1_dram_ck		,	//DDR3������ţ�ʱ����
	output									mcb1_dram_ck_n		,	//DDR3������ţ�ʱ�Ӹ�
	//  ===============================================================================================
	//  �������֣������ӿ��ź�
	//  ===============================================================================================
	input									i_flash_hold		,	//�����hold�ź�
	output									o_flash_hold		,	//�����hold�ź�
	output									o_usb_int			,	//������ţ����ӵ�3014����3014���ж��źţ��ߵ�ƽ��Ч��>100ns��clk_pixʱ����
//	output		[3:0]						ov_test				,	//������ţ�PCB���к��㣬���Թܽ�
	output									o_unused_pin		,	//ԭ��ͼ��û�з�Ƶ���ţ�sensor�ϵĸ���������Ҫ���������
	//i2c����
	inout									scl					,	//i2cʱ����
	inout									sda						//i2c������
	);

	//	ref signals

	//  ===============================================================================================
	//	-- ref ���ز�������
	//	----��Ϊlocalparam�Ĳ�������FPGA�ڲ��߼��̶��ģ���������ˣ��Ͳ�������
	//  ===============================================================================================

	//	-------------------------------------------------------------------------------------
	//	---- ref clock_reset
	//	-------------------------------------------------------------------------------------
	localparam		OSC_BUFG_CLK_PERIOD_NS		= 25	;	//osc_bufg_clk ��ʱ������

	//	-------------------------------------------------------------------------------------
	//	---- ref ctrl_channel �ڲ�����
	//	-------------------------------------------------------------------------------------
	//	-------------------------------------------------------------------------------------
	//	�̶�λ��궨��
	//	-------------------------------------------------------------------------------------
	localparam		DATA_WD_128					= 128	;	//�����������λ��128��
	localparam		DATA_WD_64					= 64	;	//�����������λ��64��
	localparam		DATA_WD_32					= 32	;	//�����������λ��32��
	localparam		SHORT_REG_WD 				= 16	;	//�̼Ĵ���λ��
	localparam		REG_WD 						= 32	;	//�Ĵ���λ��
	localparam		LONG_REG_WD 				= 64	;	//���Ĵ���λ��

	localparam		FVAL_TS_STABLE_NS			= OSC_BUFG_CLK_PERIOD_NS*3+20	;	//ʱ���ģ���fval���ص�����ģ�����ȶ�������ʱ�����ʱ��

	//	-------------------------------------------------------------------------------------
	//	I2C��������صĺ궨��
	//	-------------------------------------------------------------------------------------
	localparam		I2C_MASTER_CLOCK_FREQ_KHZ	= PIX_CLK_FREQ_KHZ	;	//i2c_topģ����ʱ��Ƶ�ʣ���λKHz
	localparam		I2C_CLOCK_FREQ_KHZ			= 400	;	//i2cʱ��Ƶ�ʣ���λKHz
	//	-------------------------------------------------------------------------------------
	//	�Ĵ���Ĭ��ֵ�궨�壬�˺궨����ֻ�ڷ���ʱ�ſ���Ϊ TRUE�����ֲ���ʱһ��ҪΪ FALSE
	//	-------------------------------------------------------------------------------------
	localparam		REG_INIT_VALUE				= "FALSE"	;	//�Ĵ�����Ĭ�ϵĳ�ʼֵ

	//	-------------------------------------------------------------------------------------
	//	---- ref io_channel parameter
	//	-------------------------------------------------------------------------------------
	//	-------------------------------------------------------------------------------------
	//	�����˲�
	//	-------------------------------------------------------------------------------------
	localparam		MAX_TRIG_FILTER_TIME_MS	= 5		;	//�����˲����ʱ�䣬��msΪ��λ
	localparam		TRIG_FILTER_WIDTH		= log2(MAX_TRIG_FILTER_TIME_MS*PIX_CLK_FREQ_KHZ+1)	;	//�����ź��˲�ģ��Ĵ������
	//	-------------------------------------------------------------------------------------
	//	������ʱ
	//	-------------------------------------------------------------------------------------
	localparam		MAX_TRIG_DELAY_TIME_MS	= 3000	;	//������ʱ���ʱ�䣬��msΪ��λ
	localparam		TRIG_DELAY_WIDTH		= log2(MAX_TRIG_DELAY_TIME_MS*PIX_CLK_FREQ_KHZ+1)		;	//�����ź���ʱģ��Ĵ������
	//	-------------------------------------------------------------------------------------
	//	ledλ�����
	//	-------------------------------------------------------------------------------------
	localparam		LED_CTRL_WIDTH			= 5     ;	//LED CTRL �Ĵ������
	//	-------------------------------------------------------------------------------------
	//	strobe_mask��ز���
	//	-------------------------------------------------------------------------------------
	localparam		STROBE_MASK_SIMULATION	= "FALSE";	//"TRUE"Ϊ����ģʽ��"FALSE"Ϊ����ģʽ
	//	-------------------------------------------------------------------------------------
	//	---- ref data_channel parameter
	//	-------------------------------------------------------------------------------------
	//	-------------------------------------------------------------------------------------
	//	���PLLʧ����ʱ�ӵ����ڣ���nsΪ��λ
	//	-------------------------------------------------------------------------------------
	localparam		PLL_CHECK_CLK_PERIOD_NS	= OSC_BUFG_CLK_PERIOD_NS	;	//pll���ʱ�ӵ�����
	//	-------------------------------------------------------------------------------------
	//	�жϵ���С���
	//	-------------------------------------------------------------------------------------
	localparam		INT_TIME_INTERVAL_MS	= 50	;	//�жϼ��
	//	-------------------------------------------------------------------------------------
	//	trigger_status=1��ʱ�䳬��1100ms��trigger_status��0
	//	��ʱʱ�����������ع�ʱ��+������ʱ��
	//	-------------------------------------------------------------------------------------
	localparam		TRIGGER_STATUS_INTERVAL=1100	;	//trigger_status=1��ʱʱ��,1100ms
	//	-------------------------------------------------------------------------------------
	//	sensor��ز������м����
	//	-------------------------------------------------------------------------------------
	localparam		SENSOR_MAX_EDGE			= (SENSOR_MAX_WIDTH>SENSOR_MAX_HEIGHT) ? SENSOR_MAX_WIDTH : SENSOR_MAX_HEIGHT;	//�ҳ��п�������һ������
	localparam		SENSOR_ALL_PIX_DIV4		= ((SENSOR_MAX_WIDTH/2)*(SENSOR_MAX_HEIGHT/2));	//Sensor��󴰿��£��������صĸ���
	//	-------------------------------------------------------------------------------------
	//	��ƽ����ز���
	//	-------------------------------------------------------------------------------------
	localparam		WB_OFFSET_WIDTH			= log2(SENSOR_MAX_EDGE+1)	;			//��ƽ��ģ��ƫ��λ�üĴ������
	localparam		WB_GAIN_WIDTH			= 11	;							//��ƽ��ģ������Ĵ������
	localparam		WB_STATIS_MAX_DIV4		= (SENSOR_ALL_PIX_DIV4*255/4);
	//�ĸ���ɫ������ÿ����ɫ���������ͳ��ֵ��ֻͳ�Ƹ�8bit�����ÿ�����ص����ֵ��255
	localparam		WB_STATIS_WIDTH			= 2+log2(WB_STATIS_MAX_DIV4+1)	;	//��ƽ��ģ��ͳ��ֵ���
	localparam		WB_RATIO				= 8		;							//��ƽ��������ӣ��˷�������Ҫ���ƶ���λ
	//	-------------------------------------------------------------------------------------
	//	�Ҷ�ͳ����ز���
	//	-------------------------------------------------------------------------------------
	localparam		GREY_OFFSET_WIDTH		= log2(SENSOR_MAX_EDGE+1)	;			//�Ҷ�ͳ��ģ��ƫ��λ�üĴ���
	localparam		GREY_STATIS_MAX_DIV4	= (SENSOR_ALL_PIX_DIV4*255);
	//�ĸ���ɫ�������������ص����ͳ��ֵ��ֻͳ�Ƹ�8bit�����ÿ�����ص����ֵ��255
	localparam		GREY_STATIS_WIDTH		= 2+log2(GREY_STATIS_MAX_DIV4+1)	;	//�Ҷ�ͳ��ģ��ͳ��ֵ���

	//	-------------------------------------------------------------------------------------
	//	---- ref frame_buffer parameter
	//	-------------------------------------------------------------------------------------
	//	-------------------------------------------------------------------------------------
	//	֡����صĺ궨��
	//	-------------------------------------------------------------------------------------
	localparam		BUF_DEPTH_WD			= 2		;	//֡�����λ��,�������֧��8֡��ȣ���һλ��λλ
//	localparam		FSIZE_WD				= 25	;	//֡��С��ȶ���
	localparam		FSIZE_WD				= 26	;	//֡��С��ȶ��� ���֧��64Mbyte��ͼ��
	localparam		BSIZE_WD				= 9		;	//һ��BURST ������ռ��λ��

	//	-------------------------------------------------------------------------------------
	//	---- ref u3_interface parameter
	//	-------------------------------------------------------------------------------------
	//	-------------------------------------------------------------------------------------
	//	u3_interface��صĺ궨��
	//	-------------------------------------------------------------------------------------
//	localparam		PACKET_SIZE_WD			= 23		;	//ͼ���Сλ��,��λ4�ֽ�
	localparam		PACKET_SIZE_WD			= 24		;	//ͼ���Сλ��,��λ4�ֽ� ���֧��64Mbyte��ͼ��
	localparam		DMA_SIZE		 		= 16'h2000	;	//DMA SIZE��С

	//	-------------------------------------------------------------------------------------
	//	ȡ��������ȡ��
	//	-------------------------------------------------------------------------------------
	function integer log2 (input integer xx);
		integer x;
		begin
			x	= xx-1 ;
			for (log2=0;x>0;log2=log2+1) begin
				x	= x >> 1;
			end
		end
	endfunction

	//  ===============================================================================================
	//	-- ref local signal defination
	//  ===============================================================================================
	//  ===============================================================================================
	//	---- ref clock reset output
	//  ===============================================================================================
	wire							w_async_rst					;	//ʱ�Ӹ�λģ��������첽��λ��ֻ�ṩ��MCB
	wire							w_sysclk_2x					;	//ʱ�Ӹ�λģ�����������ʱ�ӣ�ֻ�ṩ��MCB
	wire							w_sysclk_2x_180				;	//ʱ�Ӹ�λģ�����������ʱ�ӣ�ֻ�ṩ��MCB
	wire							w_pll_ce_0					;	//ʱ�Ӹ�λģ�����������Ƭѡ��ֻ�ṩ��MCB
	wire							w_pll_ce_90					;	//ʱ�Ӹ�λģ�����������Ƭѡ��ֻ�ṩ��MCB
	wire							w_mcb_drp_clk				;	//ʱ�Ӹ�λģ�������calib�߼�ʱ�ӣ�ֻ�ṩ��MCB
	wire							w_bufpll_mcb_lock			;	//ʱ�Ӹ�λģ�������bufpll_mcb �����źţ�ֻ�ṩ��MCB
	wire							clk_osc_bufg				;	//ʱ�Ӹ�λģ�������40MHzʱ�ӣ�ȫ�ֻ�������
	wire							reset_osc_bufg				;	//ʱ�Ӹ�λģ�������40MHzʱ�ӵĸ�λ�ź�
	wire							clk_pix						;	//ʱ�Ӹ�λģ���������������ʱ�ӣ�55Mhz
	wire							reset_pix					;	//ʱ�Ӹ�λģ���������������ʱ�ӵĸ�λ�ź�
	wire							clk_pix_2x					;	//ʱ�Ӹ�λģ���������������ʱ�ӣ�110Mhz
	wire							reset_pix_2x				;	//ʱ�Ӹ�λģ���������������ʱ�ӵĸ�λ�ź�
	wire							clk_frame_buf				;	//ʱ�Ӹ�λģ�������֡��ʱ�ӣ���gpifʱ����ͬһ��Դͷ��Ϊ�˱�֤ģ������ԣ�֡�滹��ʹ�õ�����ʱ������
	wire							reset_frame_buf				;	//ʱ�Ӹ�λģ�������֡��ʱ�ӵĸ�λ�źţ���gpifʱ����ĸ�λ�ź���ͬһ��Դͷ
	wire							clk_gpif					;	//ʱ�Ӹ�λģ�������gpif ʱ�ӣ�100MHz
	wire							reset_gpif					;	//ʱ�Ӹ�λģ�������gpif ʱ�ӵĸ�λ�ź�
	wire							reset_u3_interface			;	//ʱ�Ӹ�λģ�������u3 interface ģ�鸴λ
	wire							w_sensor_reset_done			;	//ʱ�Ӹ�λģ�������clk_osc_bufgʱ����sensor��λ����źţ����̼���ѯ���̼���ѯ���ñ�־���ܸ�λ
	//  ===============================================================================================
	//	---- ref ctrl_channel output
	//  ===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	SPI ��̬
	//	-------------------------------------------------------------------------------------
	wire							w_spi_miso_data				;	//����ͨ�������spi_sampleʱ����spi����ź�
	wire							w_spi_miso_data_en			;	//����ͨ�������spi_sampleʱ����spi����ź�ʹ���źţ���ʹ���ź�Ϊ0ʱ��miso���Ÿ���

	//	-------------------------------------------------------------------------------------
	//	I2C ����ź�
	//	-------------------------------------------------------------------------------------
	wire							w_scl_pad_i					;	//����ͨ�����룬 i2c scl ���������ź�
	wire							w_sda_pad_i					;	//����ͨ�����룬 i2c sda ���������ź�
	wire							w_scl_pad_o					;	//����ͨ�������clk_pixʱ���� i2c scl ��������ź�
	wire							w_sda_pad_o					;	//����ͨ�������clk_pixʱ���� i2c sda ��������ź�
	wire							w_scl_padoen_o				;	//����ͨ�������clk_pixʱ���� i2c scl �������ʹ��
	wire							w_sda_padoen_o				;	//����ͨ�������clk_pixʱ���� i2c sda �������ʹ��
	wire							w_i2c_ena					;	//����ͨ�������clk_pixʱ����i2c ʹ���ź�
	wire							w_trigger_start				;	//����ͨ�������clk_pixʱ����i2c������ʼ�����

	//  -------------------------------------------------------------------------------------
	//	ͨ��
	//  -------------------------------------------------------------------------------------
	wire							w_stream_enable_pix			;	//����ͨ�������clk_pixʱ�����������źţ�û����Чʱ��
	wire							w_acquisition_start_pix		;	//����ͨ�������clk_pixʱ���򣬿����źţ�û����Чʱ��
	wire							w_stream_enable_frame_buf	;	//����ͨ�������clk_frame_bufʱ�����������źţ�û����Чʱ��
	wire							w_stream_enable_gpif		;	//����ͨ�������clk_gpifʱ�����������źţ�û����Чʱ��
	//  -------------------------------------------------------------------------------------
	//	����� clk reset top
	//  -------------------------------------------------------------------------------------
	wire							w_reset_sensor				;	//����ͨ�������clk_osc_bufgʱ���򣬸�λsensorʹ���źţ�1��ʱ�����ڿ��
	//  -------------------------------------------------------------------------------------
	//	����� io channel
	//  -------------------------------------------------------------------------------------
	wire							w_trigger_mode				;	//����ͨ·�����clk_pixʱ���򣬴���ģʽ�Ĵ�����û����Чʱ������
	wire	[3:0]					wv_trigger_source			;	//����ͨ·�����clk_pixʱ���򣬴���Դ�Ĵ�����û����Чʱ������
	wire							w_trigger_soft				;	//����ͨ·�����clk_pixʱ���������Ĵ���������ͨ�������㣬�����1��ʱ������
	wire							w_trigger_active			;	//����ͨ·�����clk_pixʱ���򣬴�����Ч�ؼĴ�����û����Чʱ������
	wire	[TRIG_FILTER_WIDTH-1:0]	wv_trigger_filter_rise		;	//����ͨ·�����clk_pixʱ���������ش����˲��Ĵ�����û����Чʱ�����ƣ�����֤������Ч
	wire	[TRIG_FILTER_WIDTH-1:0]	wv_trigger_filter_fall		;	//����ͨ·�����clk_pixʱ�����½��ش����˲��Ĵ�����û����Чʱ�����ƣ�����֤������Ч
	wire	[TRIG_DELAY_WIDTH-1:0]	wv_trigger_delay			;	//����ͨ·�����clk_pixʱ���򣬴����ӳټĴ�����û����Чʱ�����ƣ�����֤������Ч
	wire	[2:0]					wv_useroutput_level			;	//����ͨ·�����clk_pixʱ�����û��Զ�������Ĵ�����û����Чʱ������
	wire							w_line2_mode				;	//����ͨ�������clk_pixʱ����line2�������ģʽ�Ĵ���
	wire							w_line3_mode				;	//����ͨ�������clk_pixʱ����line3�������ģʽ�Ĵ���
	wire							w_line0_invert				;	//����ͨ�������clk_pixʱ����line0���ԼĴ���
	wire							w_line1_invert				;	//����ͨ�������clk_pixʱ����line1���ԼĴ���
	wire							w_line2_invert				;	//����ͨ�������clk_pixʱ����line2���ԼĴ���
	wire							w_line3_invert				;	//����ͨ�������clk_pixʱ����line3���ԼĴ���
	wire	[2:0]					wv_line_source1				;	//����ͨ�������clk_pixʱ����line1�����Դѡ��Ĵ���
	wire	[2:0]					wv_line_source2				;	//����ͨ�������clk_pixʱ����line2�����Դѡ��Ĵ���
	wire	[2:0]					wv_line_source3				;	//����ͨ�������clk_pixʱ����line3�����Դѡ��Ĵ���
	wire	[4:0]					wv_led_ctrl					;	//����ͨ�������clk_pixʱ����˫ɫ�ƿ��ƼĴ���

	//  -------------------------------------------------------------------------------------
	//	����� data channel
	//  -------------------------------------------------------------------------------------
	wire							w_sensor_init_done			;	//����ͨ·�����clk_osc_bufgʱ����sensor�Ĵ�����ʼ�����
	wire	[REG_WD-1:0]			wv_pixel_format				;	//����ͨ�������clk_pixʱ���򣬿���ͨ·��������ظ�ʽ�Ĵ�����û����Чʱ�����ƣ�0x01080001:Mono8��0x01100003:Mono10��0x01080008:BayerGR8��0x0110000C:BayerGR10
	wire							w_encrypt_state				;	//����ͨ�������clk_dnaʱ���򣬼���״̬���ϵ�󱣳ֲ��䣬������Ϊ����
	wire							w_pulse_filter_en			;	//����ͨ·�����clk_pixʱ���򣬻���У���Ĵ�����û����Чʱ������
	wire	[2:0]					wv_test_image_sel			;	//����ͨ·�����clk_pixʱ���򣬲���ͼѡ��Ĵ�����û����Чʱ�����ƣ�000:��ʵͼ,001:����ͼ��1�Ҷ�ֵ֡����,110:����ͼ��2��ֹ��б����,010:����ͼ��3������б����
	wire	[1:0]					wv_interrupt_en				;	//����ͨ·�����clk_pixʱ�����ж�ʹ�ܼĴ�����û����Чʱ������
	wire	[1:0]					wv_interrupt_clear			;	//����ͨ·�����clk_pixʱ�����ж�����Ĵ�����������Ч
	wire	[WB_OFFSET_WIDTH-1:0]	wv_wb_offset_x_start		;	//����ͨ·�����clk_pixʱ���򣬰�ƽ�������Ĵ�����û����Чʱ������
	wire	[WB_OFFSET_WIDTH-1:0]	wv_wb_offset_width			;	//����ͨ·�����clk_pixʱ���򣬰�ƽ���ȼĴ�����û����Чʱ������
	wire	[WB_OFFSET_WIDTH-1:0]	wv_wb_offset_y_start		;	//����ͨ·�����clk_pixʱ���򣬰�ƽ��������Ĵ�����û����Чʱ������
	wire	[WB_OFFSET_WIDTH-1:0]	wv_wb_offset_height			;	//����ͨ·�����clk_pixʱ���򣬰�ƽ��߶ȼĴ�����û����Чʱ������
	wire	[WB_GAIN_WIDTH-1:0]		wv_wb_gain_r				;	//����ͨ·�����clk_pixʱ���򣬰�ƽ����������Ĵ�����û����Чʱ������
	wire	[WB_GAIN_WIDTH-1:0]		wv_wb_gain_g				;	//����ͨ·�����clk_pixʱ���򣬰�ƽ���̷�������Ĵ�����û����Чʱ������
	wire	[WB_GAIN_WIDTH-1:0]		wv_wb_gain_b				;	//����ͨ·�����clk_pixʱ���򣬰�ƽ������������Ĵ�����û����Чʱ������
	wire	[GREY_OFFSET_WIDTH-1:0]	wv_grey_offset_x_start		;	//����ͨ·�����clk_pixʱ���򣬻Ҷ�ֵͳ�����������Ĵ�����û����Чʱ������
	wire	[GREY_OFFSET_WIDTH-1:0]	wv_grey_offset_width		;	//����ͨ·�����clk_pixʱ���򣬻Ҷ�ֵͳ�������ȼĴ�����û����Чʱ������
	wire	[GREY_OFFSET_WIDTH-1:0]	wv_grey_offset_y_start		;	//����ͨ·�����clk_pixʱ���򣬻Ҷ�ֵͳ������������Ĵ�����û����Чʱ������
	wire	[GREY_OFFSET_WIDTH-1:0]	wv_grey_offset_height		;	//����ͨ·�����clk_pixʱ���򣬻Ҷ�ֵͳ������߶ȼĴ�����û����Чʱ������
	wire	[REG_WD-1:0]			wv_trigger_interval			;	//����ͨ·�����clk_pixʱ���򣬴����������λus,������Ч
	//  -------------------------------------------------------------------------------------
	//	����� u3v format
	//  -------------------------------------------------------------------------------------
	wire							w_chunk_mode_active_pix		;	//����ͨ·�����clk_pixʱ����chunk���ؼĴ�����û����Чʱ������
	wire							w_chunkid_en_ts				;	//����ͨ·�����clk_pixʱ����ʱ������ؼĴ�����û����Чʱ������
	wire							w_chunkid_en_fid			;	//����ͨ·�����clk_pixʱ����frame id���ؼĴ�����û����Чʱ������
	wire	[REG_WD-1:0]			wv_chunk_size_img			;	//����ͨ·�����clk_pixʱ����chunk image��С��û����Чʱ������
	wire	[REG_WD-1:0]			wv_payload_size_pix			;	//����ͨ�������clk_pixʱ�������ݵĴ�С��������ͷ��β����Э��Ҫ��64bit������ֻ����32bit���ɣ���32bit��0
	wire	[SHORT_REG_WD-1:0]		wv_roi_offset_x				;	//����ͨ�������clk_pixʱ����ͷ���е�ˮƽƫ��
	wire	[SHORT_REG_WD-1:0]		wv_roi_offset_y				;	//����ͨ�������clk_pixʱ����ͷ���еĴ�ֱƫ��
	wire	[SHORT_REG_WD-1:0]		wv_roi_pic_width			;	//����ͨ�������clk_pixʱ����ͷ���еĴ��ڿ��
	wire	[SHORT_REG_WD-1:0]		wv_roi_pic_height			;	//����ͨ�������clk_pixʱ����ͷ���еĴ��ڸ߶�
	wire	[LONG_REG_WD-1:0]		wv_timestamp_u3				;	//����ͨ�������clk_osc_bufgʱ�����ڳ��ź�����������ʱ������������4��clk_osc_bufgʱ������ȶ�����pixʱ���������8��ʱ��֮������ȶ�
	//  -------------------------------------------------------------------------------------
	//	����� frame buffer
	//  -------------------------------------------------------------------------------------
	wire	[BUF_DEPTH_WD-1:0]		wv_frame_buffer_depth			;	//����ͨ�������֡����ȣ�2-8
	wire	[REG_WD-1:0]			wv_payload_size_frame_buf		;	//����ͨ�������clk_frame_bufʱ�������ݵĴ�С��������ͷ��β����Э��Ҫ��64bit������ֻ����32bit���ɣ���32bit��0
	wire							w_chunk_mode_active_frame_buf	;	//����ͨ�������clk_frame_bufʱ����chunk���ؼĴ���
	//  -------------------------------------------------------------------------------------
	//	����� u3 interface
	//  -------------------------------------------------------------------------------------
	wire	[REG_WD-1:0]			wv_si_payload_transfer_size	;	//����ͨ·�����clk_gpifʱ���򣬵������ݿ��С,����ͨ�������δ����Чʱ������
	wire	[REG_WD-1:0]			wv_si_payload_transfer_count;	//����ͨ·�����clk_gpifʱ���򣬵������ݿ����,����ͨ�������δ����Чʱ������
	wire	[REG_WD-1:0]			wv_si_payload_final_transfer1_size	;	//����ͨ·�����clk_gpifʱ����transfer1��С,����ͨ�������δ����Чʱ������
	wire	[REG_WD-1:0]			wv_si_payload_final_transfer2_size	;	//����ͨ·�����clk_gpifʱ����transfer2��С,����ͨ�������δ����Чʱ������
	wire	[REG_WD-1:0]			wv_payload_size_gpif		;	//����ͨ�������clk_gpifʱ�������ݵĴ�С��������ͷ��β����Э��Ҫ��64bit������ֻ����32bit���ɣ���32bit��0
	wire							w_chunk_mode_active_gpif	;	//����ͨ�������clk_gpifʱ����chunk���ؼĴ���
	//  ===============================================================================================
	//  ---- ref io_channel output
	//  ===============================================================================================
	wire	[3:0]					wv_line_status				;	//����ͨ�������clk_pixʱ����line״̬�Ĵ�����IOͨ�������ָʾIO����ѡ���״̬
	wire							w_trigger					;	//����ͨ�������clk_pixʱ���򣬴����ź�

	//  ===============================================================================================
	//  ---- ref data_channel output
	//  ===============================================================================================
	wire							w_fval_data_channel			;	//����ͨ·�����clk_pixʱ���򣬳���Ч�źţ�fval���ź��Ǿ�������ͨ���ӿ���ĳ��źţ���ͷ�������leader����������Ч��ͼ�����ݣ�ͣ���ڼ䱣�ֵ͵�ƽ
	wire							w_dvalid_data_channel		;	//����ͨ·�����clk_pixʱ����������Ч�źţ���־32λ����Ϊ��Ч����
	wire	[DATA_WD_128-1:0]		wv_pix_data_data_channel	;	//����ͨ·�����clk_pixʱ����32bit���ݣ���������Ч���룬������ʱ�Ӷ���
	wire							w_fval_deser				;	//����ͨ·������⴮PLLʱ����hispi����ĳ��ź�
	wire							w_lval_deser            	;	//����ͨ·������⴮PLLʱ����hispi��������ź�
	wire							w_trigger_mode_data_mask	;	//����ͨ·������⴮PLLʱ����data_masktrigger_mode�ź�
	wire							w_trigger_status			;	//����ͨ·������⴮PLLʱ����1-�д����ź��Ҵ���֡δ�����ϣ�0-�޴����źŻ򴥷�֡������
	wire							w_deser_pll_lock			;	//����ͨ·������⴮ģ��pll_lock
	wire							w_bitslip_done				;	//����ͨ·������⴮ģ�鲢��ʱ��ʱ���򣬱߽������źţ�Ϊ1ʱ���ܿ�ʼͼ��ɼ�
	wire							w_full_frame_state			;	//����ͨ·�����clk_pixʱ��������֡״̬�źţ����̼���ѯ
	wire	[REG_WD-1:0]			wv_pixel_format_data_channel;	//����ͨ·�����clk_pixʱ����Ŀ�����ú�ģ��������ͨ�������ظ�ʽ����һ��
	wire	[WB_STATIS_WIDTH-1:0]	wv_wb_statis_r				;	//����ͨ·�����clk_pixʱ���򣬰�ƽ�������Ҷ�ֵͳ�ƼĴ�����������Чʱ������
	wire	[WB_STATIS_WIDTH-1:0]	wv_wb_statis_g				;	//����ͨ·�����clk_pixʱ���򣬰�ƽ���̷����Ҷ�ֵͳ�ƼĴ�����������Чʱ������
	wire	[WB_STATIS_WIDTH-1:0]	wv_wb_statis_b				;	//����ͨ·�����clk_pixʱ���򣬰�ƽ���������Ҷ�ֵͳ�ƼĴ�����������Чʱ������
	wire	[WB_OFFSET_WIDTH-1:0]	wv_wb_offset_width_valid	;	//����ͨ·�����clk_pixʱ���򣬰�ƽ���ȼĴ��������ƽ��ͳ��ֵͬ��һ֡ͼ��
	wire	[WB_OFFSET_WIDTH-1:0]	wv_wb_offset_height_valid	;	//����ͨ·�����clk_pixʱ���򣬰�ƽ��߶ȼĴ��������ƽ��ͳ��ֵͬ��һ֡ͼ��
	wire	[GREY_OFFSET_WIDTH-1:0]	wv_grey_offset_width_valid	;	//����ͨ·�����clk_pixʱ���򣬻Ҷ�ֵͳ�������ȼĴ�������Ҷ�ͳ��ֵͬ��һ֡
	wire	[GREY_OFFSET_WIDTH-1:0]	wv_grey_offset_height_valid	;	//����ͨ·�����clk_pixʱ���򣬻Ҷ�ֵͳ������߶ȼĴ�������Ҷ�ͳ��ֵͬ��һ֡
	wire	[GREY_STATIS_WIDTH-1:0]	wv_grey_statis_sum			;	//����ͨ·�����clk_pixʱ���򣬵ĻҶ�ֵͳ�ƼĴ�������Ҷ�ͳ��ֵ����ͬ��һ֡��������ظ�ʽΪ8bit����ֵΪ����8bitͳ��ֵ��������ظ�ʽΪ10bit����ֵΪ����10bitͳ��ֵ��
	wire	[1:0]					wv_interrupt_state			;	//����ͨ·�����clk_pixʱ�����ж�״̬�Ĵ���
	wire							w_sync_buffer_error				;	//����ͨ·�����sync_bufferģ������������ţ�����ͬ��phy��������lval��ͬʱ��������1
	//  ===============================================================================================
	//  ---- ref freq_change
	//  ===============================================================================================
	wire									w_fval_fix		;
	wire									w_data_valid_fix		;
	wire	[DATA_WD_64-1:0]				wv_pix_data_fix		;
	//  ===============================================================================================
	//  ---- ref u3v_format output
	//  ===============================================================================================
	wire									w_u3v_format_fval					;	//u3v_formatģ�������clk_pixʱ���򣬳���Ч�ź�
	wire									w_u3v_format_dvalid					;	//u3v_formatģ�������clk_pixʱ����������Ч�ź�
	wire	[DATA_WD_64-1		:0]			wv_u3v_format_data					;	//u3v_formatģ�������clk_pixʱ��������
	wire									w_trailer_flag						;	//u3v_formatģ�������clk_pixʱ����β���ź�
	//  ===============================================================================================
	//  ---- ref frame_buffer output
	//  ===============================================================================================
	wire	[DATA_WD_32-1:0]		wv_frame_buffer_data		;	//frame_bufferģ�������clk_frame_bufʱ����֡���FIFO������������32bit
	wire							w_frame_buffer_dvalid		;	//frame_bufferģ�������clk_frame_bufʱ����֡�����������Ч
	wire							w_ddr_init_done				;	//frame_bufferģ�������mcb_drp_clkʱ����MCB����ĳ�ʼ�������ź�
	wire							w_wr_error					;	//frame_bufferģ�������ʱ����δ֪����MCBӲ�������DDR�����ź�
	wire							w_rd_error					;	//frame_bufferģ�������ʱ����δ֪����MCBӲ�������DDR�����ź�
	wire							w_back_buf_empty			;	//frame_bufferģ�������clk_gpifʱ����֡����FIFO�ձ�־������ָʾ֡�����Ƿ������ݿɶ�
	wire							w_frame_buffer_fifo_full	;	//frame_bufferģ�������clk_pixʱ����֡��ǰ��FIFO ��
	wire							w_frame_buffer_front_fifo_overflow;//frame_bufferģ�������clk_pixʱ����,֡��ǰ��FIFO��� 0:֡��ǰ��FIFOû����� 1:֡��ǰ��FIFO���ֹ����������
	//  ===============================================================================================
	//  ---- ref u3_interface output
	//  ===============================================================================================
	wire									w_buf_rd							;	//u3_interfaceģ�������clk_gpifʱ���򣬶�ȡ֡����FIFO�źţ���i_data_valid�źŹ�ָͬʾ������Ч
	wire									w_usb_wr_for_led					;	//GPIF д�ź� - ��led_ctrlģ��
	wire									w_usb_pktend_n_for_test				;	//GPIF �������źţ��������������

	//  ===============================================================================================
	//  ---- ref others
	//  ===============================================================================================
	wire							w_ddr_error					;	//frame_bufferģ�������ʱ����δ֪����MCBӲ����أ�DDR�����ź�
	wire	[4:0]					wv_gpif_state				;	//GPIF ״̬
	wire	[3:0]					wv_fval_state				;	//fval ״̬


	//  ===============================================================================================
	//  ---- ref test signals
	//  ===============================================================================================


	//	ref ARCHITECTURE
	//  ===============================================================================================
	//	ref io logic
	//  ===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	flash��hold����ܽű�����holdֱ�����1
	//	-------------------------------------------------------------------------------------
	//	assign	o_flash_hold	= i_flash_hold;
	assign	o_flash_hold		= 1'b1;
	//	-------------------------------------------------------------------------------------
	//	spi ��˫������ڶ���ʵ��
	//	-------------------------------------------------------------------------------------
	assign	o_usb_spi_miso		= w_spi_miso_data_en ? w_spi_miso_data : 1'bz;

	//	-------------------------------------------------------------------------------------
	//	1.sensor��һЩ����ܽ��� 1��2 ����fpga��ֻ���õ�1����Ϊ�˵�·���ź������Կ��ǣ���һ��Ҳ��Ҫ�����������ţ���˾ͱ�����һ���߼�
	//	2.flash��hold����ܽţ�����
	//	-------------------------------------------------------------------------------------
	assign	o_unused_pin		= w_frame_buffer_fifo_full;

	//	-------------------------------------------------------------------------------------
	//	���Թܽ�
	//	-------------------------------------------------------------------------------------
//	assign	ov_test[0]		= 0;
//	assign	ov_test[1]		= 0;
//	assign	ov_test[2]		= 0;
//	assign	ov_test[3]		= 0;

	//  ===============================================================================================
	//	ref internal logic for test
	//  ===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	ddr�Ĵ���ָʾ�ź�
	//	-------------------------------------------------------------------------------------
	assign	w_ddr_error			= w_wr_error | w_rd_error;

	//	-------------------------------------------------------------------------------------
	//	gpif�ӿڵ�״̬������ʹ��
	//	-------------------------------------------------------------------------------------
	assign	wv_gpif_state[4:0]	= {2'b00,w_usb_pktend_n_for_test,w_usb_wr_for_led,i_usb_flagb_n};

	//	-------------------------------------------------------------------------------------
	//	fval state������ʹ��
	//	-------------------------------------------------------------------------------------
	assign	wv_fval_state[3:0]	= {w_back_buf_empty,w_u3v_format_fval,w_fval_data_channel,w_fval_deser};

	//	-------------------------------------------------------------------------------------
	//	i2c������̬����
	//	-------------------------------------------------------------------------------------
	assign scl	= w_i2c_ena ? (w_scl_padoen_o ? 1'bz : w_scl_pad_o) : 1'bz;
	assign sda	= w_i2c_ena ? (w_sda_padoen_o ? 1'bz : w_sda_pad_o) : 1'bz;
	assign w_scl_pad_i	= scl;
	assign w_sda_pad_i	= sda;

	assign	o_trigger	= 1'b0;

//	assign scl	= 1'bz;
//	assign sda	= 1'bz;
//	assign w_scl_pad_i	= 1'b1;
//	assign w_sda_pad_i	= 1'b1;


	//  ===============================================================================================
	//  clock_reset����
	//  ===============================================================================================
	clock_reset # (
	.DDR3_MEMCLK_FREQ		(DDR3_MEMCLK_FREQ		)
	)
	clock_reset_inst (
	//	-------------------------------------------------------------------------------------
	//	�ⲿ��������ʱ�ӣ�40MHz
	//	-------------------------------------------------------------------------------------
	.clk_osc				(clk_osc				),
	.i_reset_sensor			(w_reset_sensor			),
	.i_stream_enable		(w_stream_enable_gpif	),
	.clk_osc_bufg			(clk_osc_bufg			),
	.reset_osc_bufg			(reset_osc_bufg			),
	//	-------------------------------------------------------------------------------------
	//	MCB���ʱ��
	//	-------------------------------------------------------------------------------------
	.async_rst				(w_async_rst			),
	.sysclk_2x				(w_sysclk_2x			),
	.sysclk_2x_180			(w_sysclk_2x_180		),
	.pll_ce_0				(w_pll_ce_0				),
	.pll_ce_90				(w_pll_ce_90			),
	.mcb_drp_clk			(w_mcb_drp_clk			),
	.bufpll_mcb_lock		(w_bufpll_mcb_lock		),
	//	-------------------------------------------------------------------------------------
	//	frame_bufferʱ�ӣ�100MHz
	//	-------------------------------------------------------------------------------------
	.clk_frame_buf			(clk_frame_buf			),
	.reset_frame_buf		(reset_frame_buf		),
	//	-------------------------------------------------------------------------------------
	//	��������ʱ�ӣ�55MHz
	//	-------------------------------------------------------------------------------------
	.clk_pix				(clk_pix				),
	.reset_pix				(reset_pix				),
	//	-------------------------------------------------------------------------------------
	//	��������ʱ�ӣ�110MHz
	//	-------------------------------------------------------------------------------------
	.clk_pix_2x				(clk_pix_2x				),
	.reset_pix_2x			(reset_pix_2x			),
	//	-------------------------------------------------------------------------------------
	//	sensorʱ�ӣ�20MHz
	//	-------------------------------------------------------------------------------------
	.o_clk_sensor			(o_clk_sensor			),
	.o_sensor_reset_n		(o_sensor_reset_n		),
	.o_sensor_reset_done	(w_sensor_reset_done	),
	//	-------------------------------------------------------------------------------------
	//	USBʱ�ӣ�100MHz
	//	-------------------------------------------------------------------------------------
	.o_clk_usb_pclk			(o_clk_usb_pclk			),
	.clk_gpif				(clk_gpif				),
	.reset_gpif				(reset_gpif				),
	.reset_u3_interface		(reset_u3_interface		)
	);

	//  ===============================================================================================
	//  ctrl_channel����
	//  ===============================================================================================
	ctrl_channel # (
	.OSC_BUFG_CLK_PERIOD_NS		(OSC_BUFG_CLK_PERIOD_NS		),
	.WB_OFFSET_WIDTH			(WB_OFFSET_WIDTH			),
	.WB_GAIN_WIDTH				(WB_GAIN_WIDTH				),
	.WB_STATIS_WIDTH			(WB_STATIS_WIDTH			),
	.GREY_OFFSET_WIDTH			(GREY_OFFSET_WIDTH			),
	.GREY_STATIS_WIDTH			(GREY_STATIS_WIDTH			),
	.TRIG_FILTER_WIDTH			(TRIG_FILTER_WIDTH			),
	.TRIG_DELAY_WIDTH			(TRIG_DELAY_WIDTH			),
	.LED_CTRL_WIDTH				(LED_CTRL_WIDTH				),
	.SHORT_REG_WD				(SHORT_REG_WD				),
	.REG_WD						(REG_WD						),
	.LONG_REG_WD				(LONG_REG_WD				),
	.BUF_DEPTH_WD				(BUF_DEPTH_WD				),
	.I2C_MASTER_CLOCK_FREQ_KHZ	(I2C_MASTER_CLOCK_FREQ_KHZ	),
	.I2C_CLOCK_FREQ_KHZ			(I2C_CLOCK_FREQ_KHZ			)
	)
	ctrl_channel_inst(
	//  ===============================================================================================
	//	�����ź�
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	spiʱ����
	//  -------------------------------------------------------------------------------------
	.i_spi_clk					(i_usb_spi_sck			),
	.i_spi_cs_n					(i_spi_cs_n_fpga		),
	.i_spi_mosi					(i_usb_spi_mosi			),
	.o_spi_miso_data			(w_spi_miso_data		),
	.o_spi_miso_data_en			(w_spi_miso_data_en		),
	//  -------------------------------------------------------------------------------------
	//	40MHzʱ��
	//  -------------------------------------------------------------------------------------
	.clk_osc_bufg				(clk_osc_bufg			),
	.reset_osc_bufg				(reset_osc_bufg			),
	//  -------------------------------------------------------------------------------------
	//	pix ʱ����
	//  -------------------------------------------------------------------------------------
	.clk_pix				    (clk_pix				),
	.reset_pix					(reset_pix				),
	.i_fval						(w_fval_data_channel	),
	//  -------------------------------------------------------------------------------------
	//	frame buf ʱ����
	//  -------------------------------------------------------------------------------------
	.clk_frame_buf			    (clk_frame_buf			),
	.reset_frame_buf			(reset_frame_buf		),
	//  -------------------------------------------------------------------------------------
	//	gpif ʱ����
	//  -------------------------------------------------------------------------------------
	.clk_gpif			        (clk_gpif				),
	.reset_gpif					(reset_gpif				),
	//  ===============================================================================================
	//	���������ǼĴ���
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	ͨ��
	//  -------------------------------------------------------------------------------------
	.o_stream_enable_pix		(w_stream_enable_pix		),
	.o_acquisition_start_pix	(w_acquisition_start_pix	),
	.o_stream_enable_frame_buf	(w_stream_enable_frame_buf	),
	.o_stream_enable_gpif		(w_stream_enable_gpif		),
	//  -------------------------------------------------------------------------------------
	//	clk reset top
	//  -------------------------------------------------------------------------------------
	.o_reset_sensor				(w_reset_sensor			),
	.i_sensor_reset_done		(w_sensor_reset_done	),
	//  -------------------------------------------------------------------------------------
	//	i2c_top
	//  -------------------------------------------------------------------------------------
	.i_scl_pad					(w_scl_pad_i			),
	.o_scl_pad					(w_scl_pad_o			),
	.o_scl_padoen				(w_scl_padoen_o			),
	.i_sda_pad					(w_sda_pad_i			),
	.o_sda_pad					(w_sda_pad_o			),
	.o_sda_padoen 				(w_sda_padoen_o			),
	.o_i2c_ena					(w_i2c_ena				),
	.i_trigger					(w_trigger  			),
	.o_trigger_start			(w_trigger_start		),
	.i_trigger_mode				(w_trigger_mode_data_mask),
	//  -------------------------------------------------------------------------------------
	//	io channel
	//  -------------------------------------------------------------------------------------
	.o_trigger_mode				(w_trigger_mode			),
	.ov_trigger_source			(wv_trigger_source		),
	.o_trigger_soft				(w_trigger_soft			),
	.o_trigger_active			(w_trigger_active		),
	.ov_trigger_filter_rise		(wv_trigger_filter_rise	),
	.ov_trigger_filter_fall		(wv_trigger_filter_fall	),
	.ov_trigger_delay			(wv_trigger_delay		),
	.ov_useroutput_level		(wv_useroutput_level	),
	.o_line2_mode				(w_line2_mode			),
	.o_line3_mode				(w_line3_mode			),
	.o_line0_invert				(w_line0_invert			),
	.o_line1_invert				(w_line1_invert			),
	.o_line2_invert				(w_line2_invert			),
	.o_line3_invert				(w_line3_invert			),
	.ov_line_source1			(wv_line_source1		),
	.ov_line_source2			(wv_line_source2		),
	.ov_line_source3			(wv_line_source3		),
	.iv_line_status				(wv_line_status			),
	.ov_led_ctrl				(wv_led_ctrl			),

	//  -------------------------------------------------------------------------------------
	//	data channel
	//  -------------------------------------------------------------------------------------
	.i_deser_pll_lock			(w_deser_pll_lock				),
	.i_bitslip_done				(w_bitslip_done					),
	.o_sensor_init_done			(w_sensor_init_done				),
	.ov_pixel_format			(wv_pixel_format				),
	.i_full_frame_state			(w_full_frame_state		    	),
	.o_encrypt_state			(w_encrypt_state				),
	.o_pulse_filter_en			(w_pulse_filter_en				),
	.ov_test_image_sel			(wv_test_image_sel		    	),
	.ov_interrupt_en			(wv_interrupt_en		    	),
	.iv_interrupt_state			(wv_interrupt_state		    	),
	.ov_interrupt_clear			(wv_interrupt_clear		    	),
	.ov_wb_offset_x_start		(wv_wb_offset_x_start	    	),
	.ov_wb_offset_width			(wv_wb_offset_width		    	),
	.ov_wb_offset_y_start		(wv_wb_offset_y_start	    	),
	.ov_wb_offset_height		(wv_wb_offset_height	    	),
	.ov_wb_gain_r				(wv_wb_gain_r			    	),
	.ov_wb_gain_g				(wv_wb_gain_g			    	),
	.ov_wb_gain_b				(wv_wb_gain_b			    	),
	.iv_wb_statis_r				(wv_wb_statis_r			    	),
	.iv_wb_statis_g				(wv_wb_statis_g			    	),
	.iv_wb_statis_b				(wv_wb_statis_b			    	),
	.iv_wb_offset_width			(wv_wb_offset_width_valid   	),
	.iv_wb_offset_height		(wv_wb_offset_height_valid  	),
	.ov_grey_offset_x_start		(wv_grey_offset_x_start	    	),
	.ov_grey_offset_width		(wv_grey_offset_width	    	),
	.ov_grey_offset_y_start		(wv_grey_offset_y_start	    	),
	.ov_grey_offset_height		(wv_grey_offset_height	    	),
	.ov_trigger_interval		(wv_trigger_interval			),
	.iv_grey_statis_sum			(wv_grey_statis_sum		    	),
	.iv_grey_offset_width		(wv_grey_offset_width_valid 	),
	.iv_grey_offset_height		(wv_grey_offset_height_valid	),
//	.i_sync_buffer_error		(w_sync_buffer_error			),	//sync buffer ����߼������⣬��ʱ�����
	.i_sync_buffer_error		(1'b0							),

	//������
	.iv_fval_state				(wv_fval_state					),
	//  -------------------------------------------------------------------------------------
	//	u3v format
	//  -------------------------------------------------------------------------------------
	.o_chunk_mode_active		(w_chunk_mode_active_pix		),
	.o_chunkid_en_ts			(w_chunkid_en_ts				),
	.o_chunkid_en_fid			(w_chunkid_en_fid				),
	.ov_chunk_size_img			(wv_chunk_size_img				),
	.ov_payload_size_pix		(wv_payload_size_pix			),
	.ov_roi_offset_x			(wv_roi_offset_x				),
	.ov_roi_offset_y			(wv_roi_offset_y				),
	.ov_roi_pic_width			(wv_roi_pic_width				),
	.ov_roi_pic_height			(wv_roi_pic_height				),
	.ov_timestamp_u3			(wv_timestamp_u3				),
	//  -------------------------------------------------------------------------------------
	//	frame buffer
	//  -------------------------------------------------------------------------------------
	.ov_payload_size_frame_buf		(wv_payload_size_frame_buf		),
	.ov_frame_buffer_depth			(wv_frame_buffer_depth			),
	.o_chunk_mode_active_frame_buf	(w_chunk_mode_active_frame_buf	),
	.i_ddr_init_done				(w_ddr_init_done				),
	.i_ddr_error					(w_ddr_error					),
	.i_frame_buffer_front_fifo_overflow (w_frame_buffer_front_fifo_overflow),
	//  -------------------------------------------------------------------------------------
	//	u3 interface
	//  -------------------------------------------------------------------------------------
	.ov_si_payload_transfer_size			(wv_si_payload_transfer_size	    	),
	.ov_si_payload_transfer_count			(wv_si_payload_transfer_count	    	),
	.ov_si_payload_final_transfer1_size		(wv_si_payload_final_transfer1_size		),
	.ov_si_payload_final_transfer2_size		(wv_si_payload_final_transfer2_size		),
	.ov_payload_size_gpif					(wv_payload_size_gpif					),
	.o_chunk_mode_active_gpif				(w_chunk_mode_active_gpif				),

	//������
	.iv_gpif_state							(wv_gpif_state							)
	);

	//  ===============================================================================================
	//  io_channel����
	//  ===============================================================================================
	io_channel # (
	.TRIG_FILTER_WIDTH		(TRIG_FILTER_WIDTH		),
	.TRIG_DELAY_WIDTH		(TRIG_DELAY_WIDTH		),
	.LED_CTRL_WIDTH			(LED_CTRL_WIDTH			),
	.PIX_CLK_FREQ_KHZ		(PIX_CLK_FREQ_KHZ		), //clk_pixʱ��Ƶ��,55000KHz
	.SHORT_LINE_LENGTH_PCK	(SHORT_LINE_LENGTH_PCK	),
	.PHY_NUM				(PHY_NUM				),
	.PHY_CH_NUM				(PHY_CH_NUM				),
	.STROBE_MASK_SIMULATION	(STROBE_MASK_SIMULATION )
	)
	io_channel_inst(
	.clk					(clk_pix					),
	.i_trigger_mode			(w_trigger_mode				),
	.i_trigger_status		(w_trigger_status			),
	.i_acquisition_start	(w_acquisition_start_pix	),
	.i_stream_enable		(w_stream_enable_pix		),
	.i_trigger_mode_data_mask(w_trigger_mode_data_mask	),
	.ov_line_status			(wv_line_status				),
	.i_line2_mode			(w_line2_mode				),
	.i_line3_mode			(w_line3_mode				),
	.i_line0_invert			(w_line0_invert				),
	.i_line1_invert			(w_line1_invert				),
	.i_line2_invert			(w_line2_invert				),
	.i_line3_invert			(w_line3_invert				),
	.iv_filter_rise			(wv_trigger_filter_rise		),
	.iv_filter_fall			(wv_trigger_filter_fall		),
	.i_trigger_soft			(w_trigger_soft				),
	.iv_trigger_source		(wv_trigger_source			),
	.i_trigger_active		(w_trigger_active			),
	.iv_trigger_delay		(wv_trigger_delay			),
	.iv_line_source1		(wv_line_source1			),
	.iv_line_source2		(wv_line_source2			),
	.iv_line_source3		(wv_line_source3			),
	.iv_useroutput_level	(wv_useroutput_level		),
	.iv_led_ctrl			(wv_led_ctrl				),
	.i_optocoupler			(i_optocoupler				),
	.iv_gpio				(iv_gpio					),
	.o_optocoupler			(o_optocoupler				),
	.ov_gpio				(ov_gpio					),
	.o_f_led_gre			(o_f_led_gre				),
	.o_f_led_red			(o_f_led_red				),
	.i_usb_slwr_n			(w_usb_wr_for_led			),
	.i_fval					(w_fval_deser		        ),//hispi_if����ĳ��źţ��⴮ʱ����110MHz
	.i_lval					(w_lval_deser				),
	.i_sensor_strobe		(i_sensor_strobe			),
	.o_trigger				(w_trigger      			),
	//  -------------------------------------------------------------------------------------
	//	strobe_mask
	//  -------------------------------------------------------------------------------------
	.i_pll_lock				(w_deser_pll_lock			),	//�⴮PLL�����ź�
	//  -------------------------------------------------------------------------------------
	//	tigger_mask
	//  -------------------------------------------------------------------------------------
	.iv_trigger_interval	(wv_trigger_interval		)
	);
	//  ===============================================================================================
	//  data_channel����
	//  ===============================================================================================
	data_channel # (
	.PLL_CHECK_CLK_PERIOD_NS	(PLL_CHECK_CLK_PERIOD_NS	),
	.SER_FIRST_BIT				(SER_FIRST_BIT				),
	.END_STYLE					(END_STYLE					),
	.SER_DATA_RATE				(SER_DATA_RATE				),
	.DESER_CLOCK_ARC			(DESER_CLOCK_ARC			),
	.DESER_WIDTH				(DESER_WIDTH				),
	.CLKIN_PERIOD_PS			(CLKIN_PERIOD_PS			),
	.DATA_DELAY_TYPE			(DATA_DELAY_TYPE			),
	.DATA_DELAY_VALUE			(DATA_DELAY_VALUE			),
	.BITSLIP_ENABLE				(BITSLIP_ENABLE				),
	.PLL_RESET_SIMULATION		(PLL_RESET_SIMULATION		),
	.PHY_NUM					(PHY_NUM					),
	.PHY_CH_NUM					(PHY_CH_NUM					),
	.DIFF_TERM					(DIFF_TERM					),
	.IOSTANDARD					(IOSTANDARD					),
	.BAYER_PATTERN				(BAYER_PATTERN				),
	.SENSOR_DAT_WIDTH			(SENSOR_DAT_WIDTH			),
	.WB_OFFSET_WIDTH			(WB_OFFSET_WIDTH			),
	.WB_GAIN_WIDTH				(WB_GAIN_WIDTH				),
	.WB_STATIS_WIDTH			(WB_STATIS_WIDTH			),
	.WB_RATIO					(WB_RATIO					),
	.GREY_OFFSET_WIDTH			(GREY_OFFSET_WIDTH			),
	.GREY_STATIS_WIDTH			(GREY_STATIS_WIDTH			),
	.SHORT_REG_WD				(SHORT_REG_WD				),
	.REG_WD						(REG_WD						),
	.DATA_WD					(DATA_WD_128				),
	.TRIGGER_STATUS_INTERVAL	(TRIGGER_STATUS_INTERVAL	),
	.PIX_CLK_FREQ_KHZ			(PIX_CLK_FREQ_KHZ			),
	.INT_TIME_INTERVAL_MS		(INT_TIME_INTERVAL_MS		),
	.SENSOR_MAX_WIDTH			(SENSOR_MAX_WIDTH			)
	)
	data_channel_inst(
	//  -------------------------------------------------------------------------------------
	//	Sensor�ӿ�
	//  -------------------------------------------------------------------------------------
	.pix_clk_p					(pix_clk_p				        ),
	.pix_clk_n					(pix_clk_n				        ),
	.iv_pix_data_p				(iv_pix_data_p			        ),
	.iv_pix_data_n				(iv_pix_data_n			        ),
	//  -------------------------------------------------------------------------------------
	//	���ʱ����
	//  -------------------------------------------------------------------------------------
	.clk_pll_check				(clk_osc_bufg					),
	//  -------------------------------------------------------------------------------------
	//	�⴮ʱ����
	//  -------------------------------------------------------------------------------------
	.o_fval_deser               (w_fval_deser                   ),
	.o_lval_deser               (w_lval_deser                   ),
	.o_trigger_mode_data_mask	(w_trigger_mode_data_mask		),
	.o_trigger_status			(w_trigger_status				),
	//  -------------------------------------------------------------------------------------
	//	����ʱ����
	//  -------------------------------------------------------------------------------------
	.clk_pix					(clk_pix						),
	.reset_pix					(reset_pix						),
	.o_fval						(w_fval_data_channel			),
	.o_pix_data_en				(w_dvalid_data_channel			),
	.ov_pix_data				(wv_pix_data_data_channel		),
	//  -------------------------------------------------------------------------------------
	//	�Ĵ�������
	//  -------------------------------------------------------------------------------------
	.i_trigger_start			(w_trigger_start				),
	.i_trigger_mode				(w_trigger_mode					),
	.o_deser_pll_lock			(w_deser_pll_lock				),
	.o_bitslip_done				(w_bitslip_done					),
	.i_sensor_init_done			(w_sensor_init_done				),
	.i_acquisition_start		(w_acquisition_start_pix		),
	.i_stream_enable			(w_stream_enable_pix			),
	.o_full_frame_state			(w_full_frame_state				),
	.i_encrypt_state			(w_encrypt_state				),
	.i_pulse_filter_en			(w_pulse_filter_en				),
	.iv_roi_pic_width			(wv_roi_pic_width				),
	.iv_test_image_sel			(wv_test_image_sel				),
	.iv_pixel_format			(wv_pixel_format				),
	.ov_pixel_format			(wv_pixel_format_data_channel	),
	.o_sync_buffer_error		(w_sync_buffer_error			),
	//  -------------------------------------------------------------------------------------
	//	�ؿ�
	//  -------------------------------------------------------------------------------------
	.iv_offset_x				(wv_roi_offset_x				),
	.iv_offset_width			(wv_roi_pic_width				),
	//  -------------------------------------------------------------------------------------
	//	��ƽ��
	//  -------------------------------------------------------------------------------------
	.iv_wb_offset_x_start		(wv_wb_offset_x_start			),
	.iv_wb_offset_width			(wv_wb_offset_width				),
	.iv_wb_offset_y_start		(wv_wb_offset_y_start			),
	.iv_wb_offset_height		(wv_wb_offset_height			),
	.iv_wb_gain_r				(wv_wb_gain_r					),
	.iv_wb_gain_g				(wv_wb_gain_g					),
	.iv_wb_gain_b				(wv_wb_gain_b					),
	.ov_wb_statis_r				(wv_wb_statis_r					),
	.ov_wb_statis_g				(wv_wb_statis_g					),
	.ov_wb_statis_b				(wv_wb_statis_b					),
	.ov_wb_offset_width			(wv_wb_offset_width_valid		),
	.ov_wb_offset_height		(wv_wb_offset_height_valid		),
	//  -------------------------------------------------------------------------------------
	//	�Ҷ�ͳ��
	//  -------------------------------------------------------------------------------------
	.iv_grey_offset_x_start		(wv_grey_offset_x_start			),
	.iv_grey_offset_width		(wv_grey_offset_width			),
	.iv_grey_offset_y_start		(wv_grey_offset_y_start			),
	.iv_grey_offset_height		(wv_grey_offset_height			),
	.ov_grey_statis_sum			(wv_grey_statis_sum				),
	.ov_grey_offset_width		(wv_grey_offset_width_valid		),
	.ov_grey_offset_height		(wv_grey_offset_height_valid	),
	//  -------------------------------------------------------------------------------------
	//	�ж�
	//  -------------------------------------------------------------------------------------
	.iv_interrupt_en			(wv_interrupt_en				),
	.iv_interrupt_clear			(wv_interrupt_clear				),
	.ov_interrupt_state			(wv_interrupt_state				),
	.o_interrupt				(o_usb_int						)
	);


	//  ===============================================================================================
	//  freq_change����
	//  ===============================================================================================
	data_fix # (
	.DATA_WD_128					(DATA_WD_128					),
	.DATA_WD_64						(DATA_WD_64						)
	)
	data_fix_inst(
	.clk_pix						(clk_pix						),
	.reset_pix						(reset_pix						),
	.i_fval							(w_fval_data_channel			),
	.i_data_valid					(w_dvalid_data_channel			),
	.iv_data						(wv_pix_data_data_channel		),
	.clk_pix_2x						(clk_pix_2x						),
	.reset_pix_2x					(reset_pix_2x					),
	.o_fval							(w_fval_fix						),
	.o_data_valid					(w_data_valid_fix				),
	.ov_data						(wv_pix_data_fix				)
	);

	//  ===============================================================================================
	//  u3v_format����
	//  ===============================================================================================
	u3v_format # (
	.PIX_CLK_FREQ_KHZ				(PIX_CLK_FREQ_KHZ*2				),
	.FVAL_TS_STABLE_NS				(FVAL_TS_STABLE_NS				),
	.DATA_WD						(DATA_WD_64						),
	.SHORT_REG_WD 					(SHORT_REG_WD 					),
	.REG_WD 						(REG_WD 						),
	.LONG_REG_WD 					(LONG_REG_WD 					)
	)
	u3v_format_inst(
	.reset							(reset_pix_2x					),
	.clk							(clk_pix_2x						),
	.i_fval							(w_fval_fix						),
	.i_data_valid					(w_data_valid_fix				),
	.iv_data						(wv_pix_data_fix				),
	.i_stream_enable				(w_stream_enable_pix			),
	.i_acquisition_start     		(w_acquisition_start_pix   		),
	.iv_pixel_format         		(wv_pixel_format_data_channel	),
	.i_chunk_mode_active     		(w_chunk_mode_active_pix   		),
	.i_chunkid_en_ts         		(w_chunkid_en_ts        		),
	.i_chunkid_en_fid        		(w_chunkid_en_fid       		),
	.iv_chunk_size_img       		(wv_chunk_size_img      		),
	.iv_timestamp					(wv_timestamp_u3				),
	.iv_offset_x					(wv_roi_offset_x				),
	.iv_offset_y					(wv_roi_offset_y				),
	.iv_size_x						(wv_roi_pic_width				),
	.iv_size_y						(wv_roi_pic_height				),
	.iv_trailer_size_y				({16'h0,wv_roi_pic_height}		),
	.o_trailer_flag					(w_trailer_flag					),
	.o_fval							(w_u3v_format_fval   			),
	.o_data_valid					(w_u3v_format_dvalid 			),
	.ov_data                 		(wv_u3v_format_data      		)
	);

	//  ===============================================================================================
	//  frame_buffer ����
	//  ===============================================================================================
	frame_buffer # (
	.BUF_DEPTH_WD					(BUF_DEPTH_WD				),
	.NUM_DQ_PINS					(NUM_DQ_PINS         		),
	.MEM_BANKADDR_WIDTH				(MEM_BANKADDR_WIDTH  		),
	.MEM_ADDR_WIDTH					(MEM_ADDR_WIDTH      		),
	.DDR3_MEMCLK_FREQ				(DDR3_MEMCLK_FREQ			),
	.MEM_ADDR_ORDER					(MEM_ADDR_ORDER				),
	.SKIP_IN_TERM_CAL				(1							),
	.DDR3_MEM_DENSITY				(DDR3_MEM_DENSITY			),
	.DDR3_TCK_SPEED					(DDR3_TCK_SPEED				),
	.DDR3_SIMULATION				(DDR3_SIMULATION			),
	.DDR3_CALIB_SOFT_IP				(DDR3_CALIB_SOFT_IP			),
	.DDR3_P0_MASK_SIZE			    (DDR3_P0_MASK_SIZE			),
	.DDR3_P1_MASK_SIZE			    (DDR3_P1_MASK_SIZE			),
	.DATA_WD						(DATA_WD_64					),
	.GPIF_DAT_WIDTH					(GPIF_DAT_WIDTH				),
	.FSIZE_WD					    (FSIZE_WD					),
	.BSIZE_WD					    (BSIZE_WD					),
	.REG_WD 						(REG_WD 					)
	)
	frame_buffer_inst(
	.clk_vin						(clk_pix_2x							),
	.i_fval							(w_u3v_format_fval   				),
	.i_dval							(w_u3v_format_dvalid 				),
	.i_trailer_flag					(w_trailer_flag						),
	.iv_image_din					(wv_u3v_format_data  				),
	.i_stream_en_clk_in				(w_stream_enable_pix				),
	.o_fifo_full					(w_frame_buffer_fifo_full			),
	.clk_vout						(clk_gpif							),
	.i_buf_rd						(w_buf_rd							),
	.o_back_buf_empty				(w_back_buf_empty					),
	.ov_frame_dout					(wv_frame_buffer_data				),
	.o_frame_valid					(w_frame_buffer_dvalid				),
	.clk_frame_buf					(clk_frame_buf						),
	.reset_frame_buf				(reset_frame_buf					),
	.o_frame_buffer_front_fifo_overflow (w_frame_buffer_front_fifo_overflow),
	.i_stream_en					(w_stream_enable_frame_buf			),
	.iv_frame_depth					(wv_frame_buffer_depth				),
	.iv_payload_size_frame_buf		(wv_payload_size_frame_buf[FSIZE_WD-1:0]	),
	.iv_payload_size_pix			(wv_payload_size_pix[FSIZE_WD-1:0]			),//���ź�û��ʹ��
	.i_chunkmodeactive				(w_chunk_mode_active_frame_buf		),
	.i_async_rst					(w_async_rst						),
	.i_sysclk_2x					(w_sysclk_2x						),
	.i_sysclk_2x_180				(w_sysclk_2x_180					),
	.i_pll_ce_0						(w_pll_ce_0							),
	.i_pll_ce_90					(w_pll_ce_90						),
	.i_mcb_drp_clk					(w_mcb_drp_clk						),
	.i_bufpll_mcb_lock				(w_bufpll_mcb_lock					),
	.o_calib_done					(w_ddr_init_done					),
	.o_wr_error						(w_wr_error							),
	.o_rd_error						(w_rd_error							),
	.mcb1_dram_dq					(mcb1_dram_dq						),
	.mcb1_dram_a         			(mcb1_dram_a         				),
	.mcb1_dram_ba        			(mcb1_dram_ba        				),
	.mcb1_dram_ras_n     			(mcb1_dram_ras_n     				),
	.mcb1_dram_cas_n     			(mcb1_dram_cas_n     				),
	.mcb1_dram_we_n      			(mcb1_dram_we_n      				),
	.mcb1_dram_odt       			(mcb1_dram_odt       				),
	.mcb1_dram_reset_n   			(mcb1_dram_reset_n   				),
	.mcb1_dram_cke       			(mcb1_dram_cke       				),
	.mcb1_dram_dm        			(mcb1_dram_dm        				),
	.mcb1_dram_udqs      			(mcb1_dram_udqs      				),
	.mcb1_dram_udqs_n    			(mcb1_dram_udqs_n    				),
	.mcb1_rzq            			(mcb1_rzq            				),
	.mcb1_dram_udm       			(mcb1_dram_udm       				),
	.mcb1_dram_dqs       			(mcb1_dram_dqs       				),
	.mcb1_dram_dqs_n     			(mcb1_dram_dqs_n     				),
	.mcb1_dram_ck        			(mcb1_dram_ck        				),
	.mcb1_dram_ck_n      			(mcb1_dram_ck_n      				)
	);

	//  ===============================================================================================
	//  u3_interface����
	//  ===============================================================================================
	u3_interface # (
	.DATA_WD      					(DATA_WD_32      					),
	.REG_WD 						(REG_WD 							),
	.DMA_SIZE						(DMA_SIZE							),
	.PACKET_SIZE_WD					(PACKET_SIZE_WD						)
	)
	u3_interface_inst(
	.clk							(clk_gpif							),
	.reset							(reset_u3_interface					),
	.i_data_valid					(w_frame_buffer_dvalid				),
	.iv_data						(wv_frame_buffer_data				),
	.i_framebuffer_empty			(w_back_buf_empty					),
	.o_fifo_rd						(w_buf_rd							),
	.iv_payload_size				(wv_payload_size_gpif				),
	.i_chunkmodeactive				(w_chunk_mode_active_gpif			),
	.iv_transfer_count				(wv_si_payload_transfer_count      	),
	.iv_transfer_size				(wv_si_payload_transfer_size      	),
	.iv_transfer1_size				(wv_si_payload_final_transfer1_size	),
	.iv_transfer2_size				(wv_si_payload_final_transfer2_size	),
	.i_usb_flagb					(i_usb_flagb_n						),
	.ov_usb_fifoaddr				(ov_usb_fifoaddr					),
	.o_usb_slwr_n					(o_usb_slwr_n						),
	.ov_usb_data					(ov_usb_data						),
	.o_usb_pktend_n					(o_usb_pktend_n						),
	.o_usb_pktend_n_for_test		(w_usb_pktend_n_for_test			),
	.o_usb_wr_for_led				(w_usb_wr_for_led					)
	);

endmodule