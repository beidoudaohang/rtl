//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : driver_ad9970
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/7/15 13:26:59	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------
`define		TESTCASE	testcase_1
module driver_ad9970 ();

	//	ref signals
	//	===============================================================================================
	//	--ref parameter
	//	===============================================================================================
	parameter	CLK_UNIT_VENDOR		= `TESTCASE.CLK_UNIT_VENDOR	;
	parameter	CLK_FREQ_MHZ		= `TESTCASE.CLK_FREQ_MHZ	;

	//	===============================================================================================
	//	--ref signal
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	����
	//	-------------------------------------------------------------------------------------
	wire	[13:0]		iv_pix_data		;
	wire				i_vd			;
	wire				i_hd			;
	wire				cli_ad9970		;

	//	-------------------------------------------------------------------------------------
	//	���
	//	-------------------------------------------------------------------------------------
	wire				o_hl		;
	wire				o_h1		;
	wire				o_h2		;
	wire				o_rg		;
	
	wire				o_tckp		;
	wire				o_tckn		;
	wire				o_dout0p	;
	wire				o_dout0n	;
	wire				o_dout1p	;
	wire				o_dout1n	;

	//	ref ARCHITECTURE

	//	-------------------------------------------------------------------------------------
	//	����
	//	-------------------------------------------------------------------------------------
	assign	iv_pix_data			= `TESTCASE.iv_pix_data_ad9970	;
	assign	i_vd				= `TESTCASE.i_vd_ad9970	;
	assign	i_hd				= `TESTCASE.i_hd_ad9970	;
	
	assign	cli_ad9970			= `TESTCASE.cli_ad9970	;

	//	-------------------------------------------------------------------------------------
	//	ad9970 bfm
	//	-------------------------------------------------------------------------------------
	bfm_ad9970 bfm_ad9970 ();

	//	-------------------------------------------------------------------------------------
	//	ad9970ģ��
	//	-------------------------------------------------------------------------------------
	ad9970_module # (
	.CLK_UNIT_VENDOR	(CLK_UNIT_VENDOR				),
	.CLK_FREQ_MHZ		(CLK_FREQ_MHZ					)
	)
	ad9970_module_inst (
	.cli				(cli_ad9970						),
	.i_vd				(i_vd							),
	.i_hd				(i_hd							),
	.i_lvds_pattern_en	(bfm_ad9970.i_lvds_pattern_en	),
	.iv_lvds_pattern	(bfm_ad9970.iv_lvds_pattern		),
	.i_sync_align_loc	(bfm_ad9970.i_sync_align_loc	),
	.iv_sync_start_loc	(bfm_ad9970.iv_sync_start_loc	),
	.iv_sync_word0		(bfm_ad9970.iv_sync_word0		),
	.iv_sync_word1		(bfm_ad9970.iv_sync_word1		),
	.iv_sync_word2		(bfm_ad9970.iv_sync_word2		),
	.iv_sync_word3		(bfm_ad9970.iv_sync_word3		),
	.iv_sync_word4		(bfm_ad9970.iv_sync_word4		),
	.iv_sync_word5		(bfm_ad9970.iv_sync_word5		),
	.iv_sync_word6		(bfm_ad9970.iv_sync_word6		),
	.iv_hblk_tog1		(bfm_ad9970.iv_hblk_tog1		),
	.iv_hblk_tog2		(bfm_ad9970.iv_hblk_tog2		),
	.i_hl_mask_pol		(bfm_ad9970.i_hl_mask_pol		),
	.i_h1_mask_pol		(bfm_ad9970.i_h1_mask_pol		),
	.i_h2_mask_pol		(bfm_ad9970.i_h2_mask_pol		),
	.iv_tclk_delay		(bfm_ad9970.iv_tclk_delay		),
	.o_hl				(o_hl							),
	.o_h1				(o_h1							),
	.o_h2				(o_h2							),
	.o_rg				(o_rg							),
	.iv_pix_data		(iv_pix_data					),
	.o_tckp				(o_tckp							),
	.o_tckn				(o_tckn							),
	.o_dout0p			(o_dout0p						),
	.o_dout0n			(o_dout0n						),
	.o_dout1p			(o_dout1p						),
	.o_dout1n			(o_dout1n						)
	);





endmodule
