//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : testcase_4
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/4/10 16:50:28	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ���ڴ�С��16x16�������ź���Ч������ģʽ�µ�����״��
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module testcase_1 ();

	//	ref signals
	//	===============================================================================================
	//	--ref parameter
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	TESTCASE
	//	-------------------------------------------------------------------------------------
	parameter	TESTCASE_NUM			= "testcase_1"			;	//����ģ����Ҫʹ���ַ���

	//	-------------------------------------------------------------------------------------
	//	monitor paramter
	//	-------------------------------------------------------------------------------------
	//	parameter	MONITOR_OUTPUT_FILE_EN			= 0						;	//�Ƿ��������ļ�
	//	parameter	MONITOR_OUTPUT_FILE_PATH		= "file/mer_file/"		;	//����������Ҫд���·��
	//	parameter	CHK_INOUT_DATA_STOP_ON_ERROR	= 0						;
	//	parameter	CHK_PULSE_WIDTH_STOP_ON_ERROR	= 0						;

	//	-------------------------------------------------------------------------------------
	//	testcase parameter
	//	-------------------------------------------------------------------------------------
	//	parameter		DDR3_MEMCLK_FREQ	= 320		;	//Memory data transfer clock frequency DDR3-640:3125 DDR3-660:3030 DDR3-720:2778 DDR3-800:2500

	//	-------------------------------------------------------------------------------------
	//	dut parameter
	//	-------------------------------------------------------------------------------------
	parameter	FIFO_WIDTH	= 4		;
	parameter	FIFO_DEPTH	= 16	;


	//	===============================================================================================
	//	--ref signal
	//	===============================================================================================


	//	-------------------------------------------------------------------------------------
	//	dut signal
	//	-------------------------------------------------------------------------------------
	parameter	CLK_PERIOD				= 25	;	//ʱ��Ƶ�ʣ�40MHz

	reg									clk			= 1'b0;
	reg									reset		= 1'b0;
	reg		[7:0]						iv_din		= 'b0;
	reg									i_wr		= 1'b0;
	reg									i_rd		= 1'b0;



	//	ref ARCHITECTURE

	//	===============================================================================================
	//	ref ***tb ��ģ�鼤��***
	//	===============================================================================================

	//	-------------------------------------------------------------------------------------
	//	--ref DUT
	//	-------------------------------------------------------------------------------------
	always	#(CLK_PERIOD/2.0)		clk		= !clk;

	initial begin
		//$display($time, "Starting the Simulation...");
		//$monitor($time, "count1 is %d,count2 is %b,count3 is %h",cnt1,cnt2,cnt3);
		reset = 1'b1;
		#200
		reset = 1'b0;
		#10000
		$stop;

	end

	initial begin
		i_wr	= 1'b1;
		#700
		i_wr	= 1'b0;
		#200
		repeat (33) begin
			#100
			i_rd	= 1'b1;
			#10
			i_rd	= 1'b0;
		end

		#200
		i_wr	= 1'b1;
		i_rd	= 1'b1;
		#10
		i_wr	= 1'b0;
		i_rd	= 1'b0;

		#200
		i_wr	= 1'b1;
		i_rd	= 1'b1;
		#10
		i_wr	= 1'b0;
		i_rd	= 1'b0;

		#200
		i_wr	= 1'b1;
		i_rd	= 1'b1;
		#10
		i_wr	= 1'b0;
		i_rd	= 1'b0;
		#200
		i_wr	= 1'b1;
		#330
		i_wr	= 1'b0;

		#200
		i_wr	= 1'b1;
		i_rd	= 1'b1;
		#10
		i_wr	= 1'b0;
		i_rd	= 1'b0;

		#200
		i_wr	= 1'b1;
		i_rd	= 1'b1;
		#10
		i_wr	= 1'b0;
		i_rd	= 1'b0;

		#200
		i_wr	= 1'b1;
		i_rd	= 1'b1;
		#10
		i_wr	= 1'b0;
		i_rd	= 1'b0;

	end

	always @ (posedge clk) begin
		//		din	<= $random();
		if(!reset) begin
			iv_din	<= iv_din + 1'b1;
		end
	end



endmodule
