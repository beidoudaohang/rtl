//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : testcase_1
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/4/10 16:50:28	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ���ڴ�С��16x16�������ź���Ч������ģʽ�µ�����״��
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module testcase_1 ();

	//	ref signals
	//	===============================================================================================
	//	--ref parameter
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	TESTCASE
	//	-------------------------------------------------------------------------------------
	parameter	TESTCASE_NUM			= "testcase_1"			;	//����ģ����Ҫʹ���ַ���

	//	-------------------------------------------------------------------------------------
	//	testcase parameter
	//	-------------------------------------------------------------------------------------
	parameter	CLK_PERIOD				= 25	;	//ʱ��Ƶ�ʣ�40MHz

	//	-------------------------------------------------------------------------------------
	//	dut parameter
	//	-------------------------------------------------------------------------------------
	parameter	UART_TYPE				= "TXRX"	;	//"TX":ONLY TX."RX":ONLY RX."TXRX" or "RXTX":BOTH RX & TX
	parameter	UART_CLK_FREQ_KHZ		= 40000		;	//ʱ��Ƶ��
	parameter	UART_BAUD_RATE			= 115200	;	//������

	//	===============================================================================================
	//	--ref signal
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	dut signal
	//	-------------------------------------------------------------------------------------
	reg						uart_clk			= 1'b0;
	reg						uart_reset			= 1'b0;
	wire					uart_rx_ser			;


	//	ref ARCHITECTURE

	//	===============================================================================================
	//	ref ***tb ��ģ�鼤��***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	--ref dut
	//	-------------------------------------------------------------------------------------
	always	#(CLK_PERIOD/2.0)	uart_clk	= !uart_clk;

	initial begin
		//$display($time, "Starting the Simulation...");
		//$monitor($time, "count1 is %d,count2 is %b,count3 is %h",cnt1,cnt2,cnt3);
		uart_reset = 1'b1;
		#200
		uart_reset = 1'b0;
		#10000
		$stop;
	end

	assign	uart_rx_ser	= harness.o_uart_tx_ser;

	//	-------------------------------------------------------------------------------------
	//	--ref bfm
	//	-------------------------------------------------------------------------------------
	initial begin
		wait(uart_reset==1'b0);
		repeat(10) @ (posedge uart_clk);
		forever begin
			harness.bfm_uart.uart_wr_1byte_random();
		end
	end

	initial begin
		wait(uart_reset==1'b0);
		repeat(10) @ (posedge uart_clk);
		harness.bfm_uart.uart_rd_always();
	end



endmodule
