//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : judge
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2013/6/3 16:18:47	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :	��дģ���ٲ��߼�
//              1)  : Ϊ�˱����дģ��ͬʱ���빤��״̬��д�����ģ��
//
//              2)  : ����ʱ��μ�֡����ģ����ϸ˵���ĵ�
//
//              3)  : ack�ź���Ч״̬Ϊ1clk�ߵ�ƽ
//
//-------------------------------------------------------------------------------------------------
//`include			"judge_def.v"
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module judge (
	input				clk			,
	input				i_wr_req	,//д�����źţ�����Ч
	input				i_rd_req	,//�������źţ�����Ч
	output				o_wr_ack	,//д�����źţ�����Ч
	output				o_rd_ack	//�������źţ�����Ч
	);

	//ref signals
	reg					wr_ack_reg = 1'b0;
	reg					rd_ack_reg = 1'b0;

	//ref ARCHITECTURE

	//  -------------------------------------------------------------------------------------
	//  ��д�����ٲ�
	//	��д�����źſ����1 clk��
	//	���������ģ��������յ������źŵ��¸����ڽ������ź�����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if((i_wr_req == 1'b1)&&(wr_ack_reg == 1'b0)) begin				//д�������ˣ��һ�û����Ӧ��д����
			wr_ack_reg	<= 1'b1;
		end
		else begin
			wr_ack_reg	<= 1'b0;
		end
	end

	always @ (posedge clk) begin
		if((i_rd_req == 1'b1)&&(rd_ack_reg == 1'b0)) begin				//�ж��������ˣ��һ�û����Ӧ��������
			if(i_wr_req == 1'b1) begin									//������д����
				if(wr_ack_reg == 1'b1) begin							//�Ѿ���Ӧ��д������ô�������������
					rd_ack_reg	<= 1'b1;
				end
				else begin											//��û����Ӧд�����������������
					rd_ack_reg	<= 1'b0;
				end
			end
			else begin												//��ʱû��д���󣬿������������
				rd_ack_reg	<= 1'b1;
			end
		end
		else begin													//û�ж���������������ź�
			rd_ack_reg	<= 1'b0;
		end
	end

	assign	o_wr_ack	= wr_ack_reg;
	assign	o_rd_ack	= rd_ack_reg;



endmodule
