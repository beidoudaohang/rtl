//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : chipscope_top
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/10/27 10:21:13	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module chipscope_top (
	input				CLK			,
	input	[34:0]		TRIG0
	);

	//	ref signals
	wire	[35:0]			CONTROL0	;

	//	ref ARCHITECTURE
	chipscope_icon_user1_1port chipscope_icon_user1_1port_inst (
	.CONTROL0	(CONTROL0	)
	);

	chipscope_ila_w35_d1k chipscope_ila_w35_d1k_inst (
	.CONTROL	(CONTROL0	),
	.CLK		(CLK		),
	.TRIG0		(TRIG0		)
	);


endmodule
