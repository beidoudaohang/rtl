//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : sensor_noise
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/4/16 13:59:24	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module sensor_noise # (
	parameter			DATA_WIDTH			= 8		,	//����λ��
	parameter			CHANNEL_NUM			= 4			//ͨ����
	)
	(
	input										clk							,	//ʱ��
	input	[15:0]								iv_line_active_pix_num		,	//�п�
	input										i_fval						,	//����Ч
	input										i_lval						,	//����Ч
	input	[DATA_WIDTH*CHANNEL_NUM-1:0]		iv_pix_data					,	//��������
	output										o_fval						,	//����Ч
	output										o_lval						,	//����Ч
	output	[DATA_WIDTH*CHANNEL_NUM-1:0]		ov_pix_data						//��������
	);

	//	ref signals
	reg		[7:0]								lfsr_reg	= 8'hab;
	wire										lfsr_seed	;
	reg		[7:0]								time_cnt	= 8'b0;
	wire										noise_en	;
	wire	[DATA_WIDTH*CHANNEL_NUM-1:0]		noise_data	;


	//	ref ARCHITECTURE

	//	-------------------------------------------------------------------------------------
	//	lfsr ���������
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		lfsr_reg	<= {lfsr_reg[6:0],lfsr_seed};
	end
	assign	lfsr_seed	= lfsr_reg[0] ^ lfsr_reg[2] ^ lfsr_reg[7];

	//	-------------------------------------------------------------------------------------
	//	ʱ�������
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!i_fval) begin
			time_cnt	<= 8'h0;
		end
		else begin
			if(i_lval) begin
				if(time_cnt==lfsr_reg) begin
					time_cnt	<= 8'h0;
				end
				else begin
					time_cnt	<= time_cnt + 1'b1;
				end
			end
		end
	end

	assign	noise_en	= (i_fval==1'b1 && i_lval==1'b1 && time_cnt==lfsr_reg) ? 1'b1 : 1'b0;
	assign	noise_data	= {{(DATA_WIDTH*CHANNEL_NUM-8){1'b0}},lfsr_reg[7:0]};
	assign	o_fval		= i_fval;
	assign	o_lval		= i_lval;
	assign	ov_pix_data	= (noise_en==1'b1) ? noise_data : iv_pix_data;



endmodule
