//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : timestamp
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/12/12 16:01:50	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module timestamp # (
	parameter		LONG_REG_WD				= 64		//���Ĵ���λ��
	)
	(
	input							clk					,	//40MHzʱ��
	input							reset				,	//40MHzʱ��
	input							i_fval				,	//clk_pixʱ���򣬳���Ч�������±�������ʱ�����ov_timestamp_u3
	output	[LONG_REG_WD-1:0]		ov_timestamp_u3		,	//clk_osc_bufgʱ����ʱ�������u3v formatģ��
	input							i_timestamp_load	,	//clk_osc_bufgʱ���򣬼�⵽�����أ�����ʱ�����ov_timestamp_reg
	output	[LONG_REG_WD-1:0]		ov_timestamp_reg		//clk_osc_bufgʱ����ʱ��������Ĵ���ģ��
	);

	//	ref signals

	reg		[LONG_REG_WD-1:0]		timestamp_cnt	= {LONG_REG_WD{1'b0}};
	reg		[LONG_REG_WD-1:0]		timestamp_reg	= {LONG_REG_WD{1'b0}};
	reg		[LONG_REG_WD-1:0]		timestamp_u3	= {LONG_REG_WD{1'b0}};


	reg		[2:0]		fval_shift	= 3'b000;
	wire				fval_rise		;
	wire				fval_fall		;

	//	ref ARCHITECTURE


	//  -------------------------------------------------------------------------------------
	//	��ʱ����������fval�������غ��½���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_shift	<= {fval_shift[1:0],i_fval};
	end
	assign	fval_rise	= (fval_shift[2:1]==2'b01) ? 1'b1 : 1'b0;
	assign	fval_fall	= (fval_shift[2:1]==2'b10) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//	�ڲ�������
	//	1.��λ�ź���DCM72 lock ����֮���������������ʱ������֮��ʱ����ŻἼ��
	//	2.ʱ����40MHz��������25ns��ʱ����ĵ�λ��ns����˼�����ÿ��Ҫ�ۼ�25(0x19)
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(reset) begin
			timestamp_cnt	<= {LONG_REG_WD{1'b0}};
		end
		else begin
			timestamp_cnt	<= timestamp_cnt + 5'h19;
		end
	end

	//  -------------------------------------------------------------------------------------
	//	timestamp_reg
	//	1.i_timestamp_load���������źţ���i_timestamp_load=1��ʱ�򣬽��ڲ����������浽�˿���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(i_timestamp_load) begin
			timestamp_reg	<= timestamp_cnt;
		end
	end
	assign	ov_timestamp_reg	= timestamp_reg;

	//  -------------------------------------------------------------------------------------
	//	timestamp_u3
	//	1.��fval������ʱ�����ڲ����������浽�˿���
	//	2.��fval�½���ʱ�����ڲ����������浽�˿���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(fval_rise) begin
			timestamp_u3	<= timestamp_cnt;
		end
		else if(fval_fall) begin
			timestamp_u3	<= timestamp_cnt;
		end
	end
	assign	ov_timestamp_u3	= timestamp_u3;





endmodule
