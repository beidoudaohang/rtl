//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : circuit_dependent
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/12/17 16:06:25	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ���·״̬��أ���Ϊio���ϵĹ���������ܻ�����������⣬�ڴ�ģ���н�������źŻ�ԭ��
//						������Ҫ��U2���ݣ�ֻ��ԭ�����źţ�����ԭ����źš�
//              1)  : line0���뷴��
//				2)  : line1�������
//              3)  : gpio���벻����
//				4)  : gpio�������
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module circuit_dependent (
	//���ӵ�IO�������
	input								i_optocoupler		,	//line0�������ź�
	input	[1:0]						iv_gpio				,	//line2 3 �������ź�
	//���ӵ�io channel�ĺ�ģ��
	output								o_optocoupler_in	,	//�� i_optocoupler ȡ��
	output	[1:0]						ov_gpio_in				//���� iv_gpio
	);

	//	ref signals



	//	ref ARCHITECTURE
	//  -------------------------------------------------------------------------------------
	//	����IO���״̬��line0������Ҫ����Line2 line3���벻����
	//  -------------------------------------------------------------------------------------
	assign	o_optocoupler_in	= !i_optocoupler;
	assign	ov_gpio_in			= iv_gpio;



endmodule
