//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : triggersource_sel
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/12/1 13:21:15	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :ѡ��������ź�
//              1)  : ��3���ⴥ��ѡ��һ������Դ����֧�ֶഥ��Դ
//
//              2)  : ������ʱ���·��������߼���·����Ϊ�����ź��Ƕ�bit�������ë�����
//
//              3)  : �����ģ�����˲�ģ�飬�����źŲ������ģ�飬���ں����ģ�����ٴ�ѡ��
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module triggersource_sel (
	//ʱ��
	input				clk					,	//ʱ��
	//�Ĵ�������
	input	[3:0]		iv_trigger_source	,	//ѡ������Դ��0001-������0010-line0��0100-line2��1000-line3
	//line�����ź�
	input	[2:0]		iv_linein			,	//line�����ź�
	output				o_linein				//��������Դѡ����źţ�3·�����źű�Ϊ1��
	);

	//	ref signals
	reg			sel_result	= 1'b0;

	//	ref ARCHITECTURE
	//  -------------------------------------------------------------------------------------
	//	1.��bit����
	//	2.����������ѡ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		case(iv_trigger_source)
			4'b0010	: sel_result	<= iv_linein[0];
			4'b0100	: sel_result	<= iv_linein[1];
			4'b1000	: sel_result	<= iv_linein[2];
			default	: sel_result	<= 1'b0;
		endcase
	end

	assign	o_linein	= sel_result;



endmodule
