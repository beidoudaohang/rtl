//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : ad_horizontal_driver
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/8/9 15:48:45	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module ad_horizontal_driver (
	input			clk				,	//8������ʱ��
	input			reset			,	//����ʱ�Ӹ�λ
	input			i_hl_mask_pol	,	//hblk��Чʱ��hl�ĵ�ƽ
	input			i_h1_mask_pol	,	//hblk��Чʱ��h1�ĵ�ƽ
	input			i_h2_mask_pol	,	//hblk��Чʱ��h2�ĵ�ƽ
	input			i_hblk_n		,	//hblk�źţ�����Ч
	output			o_hl			,	//hl
	output			o_h1			,	//h1
	output			o_h2			,	//h2
	output			o_rg				//rg
	);

	//	ref signals
	reg		[2:0]		ser_cnt		= 3'b0;
	reg					hl_reg		= 1'b0;
	reg					h1_reg		= 1'b0;
	reg					h2_reg		= 1'b0;

	//	ref ARCHITECTURE

	//	-------------------------------------------------------------------------------------
	//	���л�������
	//	1.ÿ��ͨ���Ĵ�������8bit����˼�������3bit����0��7�ۼ�
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(reset) begin
			ser_cnt	<= 3'b0;
		end
		else begin
			ser_cnt	<= ser_cnt + 1'b1;
		end
	end

	//	-------------------------------------------------------------------------------------
	//	hl
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(i_hblk_n==1'b0) begin
			hl_reg	<= i_hl_mask_pol;
		end
		else begin
			if(ser_cnt==3'd1) begin
				hl_reg	<= 1'b0;
			end
			else if(ser_cnt==3'd5) begin
				hl_reg	<= 1'b1;
			end
		end
	end
	assign	o_hl	= hl_reg;
	assign	o_rg	= !hl_reg;
	
	//	-------------------------------------------------------------------------------------
	//	h1
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(i_hblk_n==1'b0) begin
			h1_reg	<= i_h1_mask_pol;
		end
		else begin
			if(ser_cnt==3'd1) begin
				h1_reg	<= 1'b0;
			end
			else if(ser_cnt==3'd5) begin
				h1_reg	<= 1'b1;
			end
		end
	end
	assign	o_h1	= h1_reg;

	//	-------------------------------------------------------------------------------------
	//	h2
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(i_hblk_n==1'b0) begin
			h2_reg	<= i_h2_mask_pol;
		end
		else begin
			if(ser_cnt==3'd1) begin
				h2_reg	<= 1'b0;
			end
			else if(ser_cnt==3'd5) begin
				h2_reg	<= 1'b1;
			end
		end
	end
	assign	o_h2	= h2_reg;

endmodule
