//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : pulse_filter_rd
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/2/11 15:44:38	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ��ģ����Ҫ�����Ǵ�bufferģ���ȡ���ݣ�������4����Ҫ�Ĳ���
//              1)  : �����߼����֣��������г��źű��ص���ȡ�������Ϳ��Ƽ�����
//
//              2)  : RAM�������֣�������RAM�ĸ�λ����ʹ�ܡ���ַ
//
//              3)  : ���ѡ�񲿷֣�ѡ�� upper line��mid line������mid line�ǽ�Ҫ���˲����С�lower line��wrģ���ṩ�ġ�
//
//				4)  : ֡β��������2�У���i_fval����ʱ����Ҫ������2��lval
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module pulse_filter_rd # (
	parameter					COMPARE_LVAL_DELAY	= 5		,	//�� compare ģ���lval����ʱ
	parameter					LINE_HIDE_PIX_NUM	= 30	,	//�������ɵ�2�У���������ֵ
	parameter					LINE2FRAME_PIX_NUM	= 10	,	//�������ɵ�2�У����һ�е��½�����o_fval���½��صľ���
	parameter					SENSOR_DAT_WIDTH	= 10	,	//sensor ���ݿ��
	parameter					SHORT_REG_WD		= 16		//�̼Ĵ���λ��
	)
	(
	input								clk					,	//����ʱ��
	input	[SHORT_REG_WD-1:0]			iv_roi_pic_width	,	//�п��
	input								i_fval				,	//���ź�
	input								i_lval				,	//���ź�
	output								o_reset_buffer		,	//ram ��λ
	output	[3:0]						ov_buffer_rd_en		,	//ram ��ʹ��
	output	[11:0]						ov_buffer_rd_addr	,	//ram ����ַ
	input	[9:0]						iv_buffer_rd_dout0	,	//ram0 �������
	input	[9:0]						iv_buffer_rd_dout1	,	//ram1 �������
	input	[9:0]						iv_buffer_rd_dout2	,	//ram2 �������
	input	[9:0]						iv_buffer_rd_dout3	,	//ram3 �������
	output								o_fval				,	//�������Ч
	output								o_lval				,	//�������Ч
	output	[SENSOR_DAT_WIDTH-1:0]		ov_upper_line		,	//����Ƚ���-�����һ��
	output	[SENSOR_DAT_WIDTH-1:0]		ov_mid_line				//����Ƚ���-�м��һ��
	);

	//	ref signals

	//	-------------------------------------------------------------------------------------
	//	���ز���
	//	1.��ģ�����ʱ������=�涨�ĵ���ʱ������+�����ģ���o_lval��ɵ���ʱ������
	//	-------------------------------------------------------------------------------------
	localparam		LINE2FRAME_PIX_NUM_RD	= (LINE2FRAME_PIX_NUM+COMPARE_LVAL_DELAY);


	reg									lval_dly0			= 1'b0;
	reg									lval_dly1			= 1'b0;
	reg									lval_dly2			= 1'b0;
	wire								lval_fall			;
	reg									lval_trailer_dly0	= 1'b0;
	reg									lval_trailer_dly1	= 1'b0;
	wire								lval_trailer_fall	;
	reg									fval_dly0			= 1'b0;
	wire								fval_fall			;
	wire								fval_extend			;
	reg									lval_reg			= 1'b0;

	reg		[1:0]						lval_cnt			= 2'b0;
	reg		[1:0]						lval_cnt_dly0		= 2'b0;
	reg		[1:0]						lval_cnt_dly1		= 2'b0;
	reg									fval_reg			= 1'b0;
	reg		[1:0]						buffer_rd_en		= 2'b0;
	reg		[11:0]						buffer_rd_addr		= 12'b0;
	reg		[9:0]						upper_line_reg		= 10'b0;
	reg		[9:0]						mid_line_reg		= 10'b0;

	reg									gen_2line			= 1'b0;
	reg		[4:0]						gen_2line_hide_cnt	= 5'b0;
	reg		[11:0]						gen_2line_valid_cnt	= 12'b0;
	reg									lval_trailer		= 1'b0;
	reg		[1:0]						lval_trailer_cnt	= 2'b0;


	//	ref ARCHITECTURE

	//  ===============================================================================================
	//	ref ***ȡ����***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	�ж�����lval�ı���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		lval_dly0	<= i_lval;
		lval_dly1	<= lval_dly0;
	end
	assign	lval_fall	= (lval_dly0==1'b1 && i_lval==1'b0) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//	�ж�����fval�ı���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_dly0	<= i_fval;
	end
	assign	fval_fall	= (fval_dly0==1'b1 && i_fval==1'b0) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//	�ж�lval_trailer�ı���
	//	1.lval_trailer����֡β�������ɵ����ź�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		lval_trailer_dly0	<= lval_trailer;
		lval_trailer_dly1	<= lval_trailer_dly0;
	end
	assign	lval_trailer_fall	= (lval_trailer_dly0==1'b1 && lval_trailer==1'b0) ? 1'b1 : 1'b0;

	//  ===============================================================================================
	//	ref ***֡β��������2��***
	//	1.rd ģ��Ὣlval�ź����ƽ��2�У��� i_fval=0ʱ��i_lvalҲΪ0��ֻ����ģ���ڲ���������2�� lval
	//	2.�Ĵ�����������Ч���������̶�Ϊ���������fval��lval�½���֮��ľ����ɲ�������
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	gen_2line ����֡β2�еı�־
	//	1.��i_fval�½���ʱ����־��λ
	//	2.���Ѿ�������2��lval����lval��fval֮��ľ����������ʱ����־����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(fval_fall) begin
			gen_2line	<= 1'b1;
		end
		else begin
			if(lval_trailer_cnt==2'b10 && gen_2line_hide_cnt==(LINE2FRAME_PIX_NUM_RD+1)) begin
				gen_2line	<= 1'b0;
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	������֡β2�е�����������
	//	1.��������־=0ʱ������������
	//	2.��������־=1�Ҳ�����lval=0ʱ������������
	//	2.��������־=1�Ҳ�����lval=1ʱ������������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!gen_2line) begin
			gen_2line_hide_cnt	<= 5'b0;
		end
		else begin
			if(!lval_trailer) begin
				gen_2line_hide_cnt	<= gen_2line_hide_cnt + 1'b1;
			end
			else begin
				gen_2line_hide_cnt	<= 5'b0;
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	������֡β2�е�����Ч������
	//	1.��������־=0ʱ������������
	//	2.��������־=1�Ҳ�����lval=0ʱ������������
	//	3.�˴������ж� gen_2line ��״̬����Ϊ�� gen_2line=0ʱ�� lval_trailer Ҳ����0
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!lval_trailer) begin
			gen_2line_valid_cnt	<= 5'b0;
		end
		else begin
			gen_2line_valid_cnt	<= gen_2line_valid_cnt + 1'b1;
		end
	end

	//  -------------------------------------------------------------------------------------
	//	�����ɵ�lval
	//	1.��������������������������ֵʱ��lval��Ϊ1
	//	2.���Ѿ�������2��lval����ôlval_trailerһ��Ҫ���0
	//	3.����û�в���2��lvalʱ��
	//	--3.1����Ч�������������п��-1ʱ��lval��Ϊ0
	//	--3.2����������if���ʽ֮�У�����������߼�·������ʡ��reg��fmax������180����
	//	4.������ж� lval cnt�������� hide cnt �� valid cnt ʱ�������������⣺
	//	--��LINE2FRAME_PIX_NUM_RD����LINE_HIDE_PIX_NUMʱ���ͻ�������1��lval����ȻĿǰ�Ĳ������������������������
	//	--����Ϊ��ģ���ͨ���Կ��ǣ�����Ӧ�ü��� lval_cnt �������ж�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!gen_2line) begin
			lval_trailer	<= 1'b0;
		end
		else begin
			if(lval_trailer_cnt==2'b10) begin
				lval_trailer	<= 1'b0;
			end
			else begin
				if(gen_2line_hide_cnt==(LINE_HIDE_PIX_NUM-1)) begin
					lval_trailer	<= 1'b1;
				end
				else if(gen_2line_valid_cnt==(iv_roi_pic_width[11:0]-1)) begin
					lval_trailer	<= 1'b0;
				end
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	lval_trailer_cnt
	//	1.�� lval_trailer ���½��ؼ���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!gen_2line) begin
			lval_trailer_cnt	<= 2'b0;
		end
		else begin
			if(lval_trailer_fall) begin
				lval_trailer_cnt	<= lval_trailer_cnt + 1'b1;
			end
		end
	end

	//  ===============================================================================================
	//	ref ***�����г��ź�***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//                  ______________________________________________________________
	//	i_fval         _|                                                            |_____________________________
	//                                                                               __________________
	//  gen_2line      ______________________________________________________________|                |____________
	//                  _______________________________________________________________________________
	//	fval_extend    _|                                                                             |____________
	//                      ____    ____      ____    ____            ____    ____
	//	i_lval         _____|  |____|  |______|  |____|  |____....____|  |____|  |_________________________________
	//                                                                                  ____    ____
	//	lval_gen       _________________________________________________________________|  |____|  |_______________
	//
	//                                    _____________________________________________________________
	//	o_fval         ___________________|                                                           |____________
	//
	//                                        ____    ____            ____    ____      ____    ____
	//	o_lval         _______________________|  |____|  |____....____|  |____|  |______|  |____|  |_______________
	//
	//  -------------------------------------------------------------------------------------
	//  -------------------------------------------------------------------------------------
	//	fval_extend - չ��֮���fval
	//	1.gen_2line����i_fval�½��ز�����
	//	2.fval_dly0 �� gen_2line �ĸߵ�ƽ֮���νӽ��ܣ�û�е͵�ƽ
	//	3.fval_extend �� i_fval ��ȣ������ʱ1�ģ�֡β�����2�е�ʱ��
	//  -------------------------------------------------------------------------------------
	assign	fval_extend		= fval_dly0 | gen_2line;

	//  -------------------------------------------------------------------------------------
	//	lval���ؼ�����
	//	1.��չ���� fval =0 ʱ��lval_cnt ����
	//	2.��չ���� fval =1 ʱ���� i_lval ���½��� ���� �������ɵ� lval_trailer ���½���ʱ������������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!fval_extend) begin
			lval_cnt	<= 2'b00;
		end
		else begin
			if(lval_fall==1'b1 || lval_trailer_fall==1'b1) begin
				lval_cnt	<= lval_cnt + 1'b1;
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	fval_reg - ����ĳ��ź�
	//	1.��i_fval=0��gen_2line=0ʱ�����ܽ�fval_reg����
	//	2.֡��Ч����֮��fval_reg=1
	//	3.o_fval �� i_fval ��ȣ����ƽ����2��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!fval_extend) begin
			fval_reg	<= 1'b0;
		end
		else if(lval_cnt==2'b10) begin
			fval_reg	<= 1'b1;
		end
	end
	assign	o_fval	= fval_reg;

	//  -------------------------------------------------------------------------------------
	//	��������lval
	//	1.��o_fval=0ʱ��o_lval=0
	//	2.�����ɵ�lval���� (1)������ǰ���е�ԭʼi_lval (2)֡β�������ɵ�����
	//	3.ram ���ź���i_lval��lval_trailer����֮����źţ�ram��ʱ1��ʱ�����ڣ�ram�����������dly1�Ƕ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!fval_reg) begin
			lval_reg	<= 1'b0;
		end
		else begin
			lval_reg	<= lval_dly1|lval_trailer_dly1;
		end
	end
	assign	o_lval	= lval_reg;

	//  -------------------------------------------------------------------------------------
	//	�ӳ� lval cnt
	//	1.ram�����1��ʱ����ʱ
	//	2.ram���źŸ��� lval_cnt�л�
	//	3.��lval�ı�ʱ��ram���źŲ��������л���Ҫ�ӳ�2��ʱ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		lval_cnt_dly0	<= lval_cnt;
		lval_cnt_dly1	<= lval_cnt_dly0;
	end

	//  ===============================================================================================
	//	ref ***RAM�Ĳ���***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	-- ref RAM ��λ
	//	1.������֡����ʱ����λRAM�� fval_extend ��ԭʼ��i_fval��2��ʱ�䣬��Ϊǰ2��ҲҪд�뵽ram�У����ܸ�λ
	//	2.��֡��Ч����һ������Ч���д�Լ10��ʱ�ӵ�ʱ�䣬��Ҫ��֤FIFO�ܹ��Ӹ�λ״̬�ָ�����
	//  -------------------------------------------------------------------------------------
	assign	o_reset_buffer	= !fval_extend;

	//  -------------------------------------------------------------------------------------
	//	-- ref RAM ��
	//	1.��֡����ʱ�����ź�ȫΪ�� ���˴���Ҫ�� o_fval��Ϊʹ�ܣ���Ϊǰ�����ǲ�����
	//	2.��֡��Чʱ������lval cntѡȡ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!fval_reg) begin
			buffer_rd_en	<= 2'b00;
		end
		else begin
			case(lval_cnt[0])
				1'b0	: buffer_rd_en	<= {1'b0,i_lval|lval_trailer};
				1'b1	: buffer_rd_en	<= {i_lval|lval_trailer,1'b0};
				default	: buffer_rd_en	<= 2'b00;
			endcase
		end
	end
	assign	ov_buffer_rd_en[0]	= buffer_rd_en[0];
	assign	ov_buffer_rd_en[2]	= buffer_rd_en[0];
	assign	ov_buffer_rd_en[1]	= buffer_rd_en[1];
	assign	ov_buffer_rd_en[3]	= buffer_rd_en[1];

	//  -------------------------------------------------------------------------------------
	//	-- ref RAM ����ַ
	//	1.��֡��Чʱ����ʹ����i_lvalʱ����������ַҪ֮��һ��ʱ���ٱ仯
	//	2.���������ɵ�2���£�ҲҪ��ram
	//	3.��֡����ʱ��ram����ַ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(fval_reg) begin
			if(lval_dly0==1'b1 || lval_trailer_dly0==1'b1) begin
				buffer_rd_addr	<= buffer_rd_addr + 1'b1;
			end
			else if(lval_dly0==1'b0 || lval_trailer_dly0==1'b0) begin
				buffer_rd_addr	<= 12'h0;
			end
		end
		else begin
			buffer_rd_addr	<= 12'h0;
		end
	end
	assign	ov_buffer_rd_addr	= buffer_rd_addr;

	//  ===============================================================================================
	//	ref ***���ѡ��***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	ѡ���������һ������
	//	1.֡��Чʱ������lval_cnt��״̬��ѡ��ram
	//	2.֡����ʱ�������������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(fval_reg) begin
			case(lval_cnt_dly1)
				2'b10	: upper_line_reg	<= iv_buffer_rd_dout2;
				2'b11	: upper_line_reg	<= iv_buffer_rd_dout3;
				2'b00	: upper_line_reg	<= iv_buffer_rd_dout0;
				2'b01	: upper_line_reg	<= iv_buffer_rd_dout1;
				default	: upper_line_reg	<= 10'b0;
			endcase
		end
		else begin
			upper_line_reg	<= 10'b0;
		end
	end
	assign	ov_upper_line	= upper_line_reg[SENSOR_DAT_WIDTH-1:0];

	//  -------------------------------------------------------------------------------------
	//	���ѡ����м�������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(fval_reg) begin
			case(lval_cnt_dly1)
				2'b10	: mid_line_reg	<= iv_buffer_rd_dout0;
				2'b11	: mid_line_reg	<= iv_buffer_rd_dout1;
				2'b00	: mid_line_reg	<= iv_buffer_rd_dout2;
				2'b01	: mid_line_reg	<= iv_buffer_rd_dout3;
				default	: mid_line_reg	<= 10'b0;
			endcase
		end
		else begin
			mid_line_reg	<= 10'b0;
		end
	end
	assign	ov_mid_line	= mid_line_reg[SENSOR_DAT_WIDTH-1:0];


endmodule
