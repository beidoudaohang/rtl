//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : ccd_sharp_vshift
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/8/10 14:14:50	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module ccd_sharp_vshift (
	input			xv1				,	//��ֱ����
	input			xv2				,	//��ֱ����
	input			xv3				,	//��ֱ����
	input			xv4				,	//��ֱ����
	input			xsg				,	//�ع�����ź�
	output			o_line_change	,	//��ֱ��ת����
	output			o_frame_change		//�ع�����ź�
	);

	//	ref signals
	wire	[3:0]		xv_comb		;
	reg					line_change		= 1'b0;
	reg					frame_change	= 1'b0;

	//	ref ARCHITECTURE

	//	-------------------------------------------------------------------------------------
	//	��ֱ��ת
	//	-------------------------------------------------------------------------------------
	assign	xv_comb	= {xv4,xv3,xv2,xv1};

	initial begin
		forever begin
			line_change	= 1'b0;
			wait(xv_comb==4'b0011);
			wait(xv_comb==4'b0111);
			wait(xv_comb==4'b0110);
			wait(xv_comb==4'b1110);
			wait(xv_comb==4'b1100);
			wait(xv_comb==4'b1101);
			wait(xv_comb==4'b1001);
			wait(xv_comb==4'b1011);
			wait(xv_comb==4'b0011);
			#10
			line_change	= 1'b1;
			#10
			line_change	= 1'b0;
		end
	end
	assign	o_line_change	= line_change;

	//	-------------------------------------------------------------------------------------
	//	�ع�
	//	-------------------------------------------------------------------------------------
	initial begin
		forever begin
			frame_change	= 1'b0;
			@(negedge xsg)
			#10
			frame_change	= 1'b1;
			#10
			frame_change	= 1'b0;
		end
	end
	assign	o_frame_change	= frame_change;


endmodule
