//-------------------------------------------------------------------------------------------------
//  -- Corporation  : MicroRTL.com
//  -- Email        : haitaox2013@gmail.com
//  -- Module       :
//-------------------------------------------------------------------------------------------------
//  -- Description  :
//
//-------------------------------------------------------------------------------------------------
//  -- Changelog    :
//  -- Author       | Date                  | Content
//  -- Michael      | 2014/12/8 14:44:37	|
//-------------------------------------------------------------------------------------------------
//`include			"_def.v"
//time unit/precision
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module uart_tx_bit (
	input				clk				,	//��ʱ�ӣ������� i_16x_baud_en ��2��
	input				i_16x_baud_en	,	//�����ʵ�16������ʹ���źţ��ߵ�ƽ��Ч��1��clk�Ŀ��
	input	[7:0]		iv_fifo_dout	,	//fifo���������
	input				i_fifo_empty	,	//fifo�Ŀ��ź�
	output				o_fifo_rd		,	//��fifo�ź�
	output				o_uart_tx_ser		//uart���Ͷ˿�
	);

	//	ref signals
	reg		[3:0]		en_16_cnt	= 4'b0;
	reg		[3:0]		tx_bit_cnt	= 4'b0;
	reg					fifo_rd_int	= 1'b0;
	reg		[9:0]		shift_reg	= 10'b0;
	reg					state_cnt	= 1'b0;

	//	ref ARCHITECTURE


	//  -------------------------------------------------------------------------------------
	//	ÿ��bit��ʱ���൱��16�� i_16x_baud_en
	//	������״̬1(��λ)ʱ���������ۼ�
	//	������״̬0(��fifo)ʱ������������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(state_cnt) begin
			if(i_16x_baud_en) begin
				en_16_cnt	<= en_16_cnt + 1'b1;
			end
		end
		else begin
			en_16_cnt	<= 'b0;
		end
	end

	//  -------------------------------------------------------------------------------------
	//	���͵� bit �ļ�����
	//	������״̬1(��λ)ʱ��ÿ����16�Σ�����һ��
	//	������״̬0(��fifo)ʱ������������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(state_cnt) begin
			if((i_16x_baud_en==1'b1)&&(en_16_cnt==4'b1111)) begin
				tx_bit_cnt	<= tx_bit_cnt + 1'b1;
			end
		end
		else begin
			tx_bit_cnt	<= 'b0;
		end
	end

	//  -------------------------------------------------------------------------------------
	//	��fifo��1��ʱ�ӿ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if((state_cnt==1'b0)&&(i_fifo_empty==1'b0)&&(i_16x_baud_en==1'b1)) begin
			fifo_rd_int	<= 1'b1;
		end
		else begin
			fifo_rd_int	<= 1'b0;
		end
	end
	assign	o_fifo_rd	= fifo_rd_int;

	//  -------------------------------------------------------------------------------------
	//	��λ�Ĵ���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(state_cnt) begin
			if((i_16x_baud_en==1'b1)&&(en_16_cnt==4'b1111)) begin
				shift_reg	<= {shift_reg[0],shift_reg[9:1]};
			end
		end
		else begin
			shift_reg	<= {1'b1,iv_fifo_dout,1'b0};	//stop + 8bit + start
		end
	end
	assign	o_uart_tx_ser	= (state_cnt==1'b1) ? shift_reg[0] : 1'b1;

	//  -------------------------------------------------------------------------------------
	//	״̬�ж�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		case(state_cnt)
			//  -------------------------------------------------------------------------------------
			//	״̬0-��fifo����״̬�൱�ڸ�λ�Ĵ�����״̬
			//  -------------------------------------------------------------------------------------
			1'b0 : begin
				if((i_fifo_empty==1'b0)&&(i_16x_baud_en==1'b1)) begin
					state_cnt	<= 1'b1;
				end
				else begin
					state_cnt	<= 1'b0;
				end
			end
			//  -------------------------------------------------------------------------------------
			//	״̬1-��λ
			//  -------------------------------------------------------------------------------------
			1'b1 : begin
				if((i_16x_baud_en==1'b1)&&(en_16_cnt==4'b1111)&&(tx_bit_cnt==4'b1001)) begin
					state_cnt	<= 1'b0;
				end
				else begin
					state_cnt	<= 1'b1;
				end
			end
			default : begin

			end
		endcase
	end

endmodule
