//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : interupt
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/12/5 15:54:33	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : �жϹ���ģ��
//              1)  : �����ж�״̬���ж�����
//
//              2)  : 3014���ж����Ÿ���Ч���ߵ�ƽ����100ns
//
//              3)  : �ж�����ʱ������֮���һ������֡������ж��ź�
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module interrupt # (
	parameter		REG_WD					= 32		,	//�Ĵ���λ��
	parameter		INT_TIME_INTERVAL_MS	= 50		,	//�жϼ��
	parameter		CLK_FREQ_KHZ			= 55000			//����ʱ��Ƶ�ʣ���λKHZ���ܶ�ģ���ø�ʱ����Ϊ��ʱ������˱���д������ʱ�ӵ�Ƶ��
	)
	(
	//Sensor�����ź�
	input					clk					,	//����ʱ��
	input					i_fval				,	//���źţ��Ҷ�ͳ��ģ�����
	//�ж���ؼĴ���
	input					i_acquisition_start	,	//�����źţ�0-ͣ�ɣ�1-����
	input					i_stream_enable		,	//��ʹ���źţ�0-ͣ�ɣ�1-����
	input					i_interrupt_en_grey	,	//2a�ж�ʹ�ܣ�����Ч
	input					i_interrupt_en_wb	,	//��ƽ���ж�ʹ�ܣ�����Ч
	input	[1:0]			iv_interrupt_clear	,	//�ж��������źţ�����Ч������ͨ�������㣬bit0-��2a�жϣ�bit1-���ƽ���ж�
	output	[1:0]			ov_interrupt_state	,	//�ж�״̬�����ж�ʹ�ܶ�Ӧ������Ч��bit0-2a�ж�״̬��bit1-��ƽ���ж�״̬
	output					o_interrupt				//�����ⲿ���ж��źţ��ж�Ƶ��20Hz���¡�����Ч�����������100ns
	);

	//	ref signals
	localparam	TIME_INTERVAL	= INT_TIME_INTERVAL_MS*CLK_FREQ_KHZ	;	//������ INT_TIME_INTERVAL_MS ����Ҫ���ٸ�ʱ������
	localparam	CNT_WIDTH		= log2(TIME_INTERVAL+1)	;	//������λ��

	//	-------------------------------------------------------------------------------------
	//	ȡ��������ȡ��
	//	-------------------------------------------------------------------------------------
	function integer log2 (input integer xx);
		integer x;
		begin
			x	= xx-1 ;
			for (log2=0;x>0;log2=log2+1) begin
				x	= x >> 1;
			end
		end
	endfunction

	reg		[1:0]				fval_shift				= 2'b0;
	wire						fval_rise				;
	wire						fval_fall				;
	reg							fval_fall_dly0			= 1'b0;
	reg							fval_fall_dly1			= 1'b0;
	reg							fval_rise_reg			= 1'b0;
	reg							full_frame_state		= 1'b0;
	reg		[1:0]				internal_state			= 2'b0;
	reg		[1:0]				interface_state			= 2'b0;
	reg		[CNT_WIDTH-1:0]		div_time_interval_cnt	= TIME_INTERVAL;
	reg							time_up					= 1'b0;
	reg							int_rise				= 1'b0;
	reg		[4:0]				extend_int_cnt			= 5'b10000;	//Ĭ��ֵ�����ֵ����֤�ж�������ϵ��ʱ���ǵ͵�ƽ
	reg							interrupt_reg			= 1'b0;

	//	ref ARCHITECTURE

	//  ===============================================================================================
	//	ref ***ȡ����***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	fval ȡ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_shift	<= {fval_shift[0],i_fval};
	end
	assign	fval_rise	= (fval_shift[1:0]==2'b01) ? 1'b1 : 1'b0;
	assign	fval_fall	= (fval_shift[1:0]==2'b10) ? 1'b1 : 1'b0;

	//	-------------------------------------------------------------------------------------
	//	fval��ʱ�ź�
	//	1.fval_fall			- fval�½��أ������ƶ�����֡״̬
	//	2.fval_fall_dly0	- fval��һ�ģ������ƶ��ڲ��ж�״̬
	//	3.fval_fall_dly1	- fval�����ģ������ƶ��ж����ŵ�״̬
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_fall_dly0	<= fval_fall;
		fval_fall_dly1	<= fval_fall_dly0;
	end

	//  ===============================================================================================
	//	ref ***����֡***
	//	1.�����������źŶ�ʹ��ʱ������һ��fval�����غ�һ��fval�½��أ�����Ϊ��1������֡
	//	2.�����Ͱѿ���֮��ĵ�һ֡���ж϶�������ʹ������֡��Ҳ�ᶪ�������Ƕ���3a��˵Ӱ�첻����Ҫ���Ǳ�֤����֡
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	fval �����ؼĴ���
	//	1.��ʹ����Чʱ���Ĵ�������
	//	2.��ʹ����Чʱ����fval�����ص�ʱ�򣬼Ĵ�����1
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if((i_acquisition_start&i_stream_enable)==1'b0) begin
			fval_rise_reg	<= 1'b0;
		end
		else begin
			if(fval_rise) begin
				fval_rise_reg	<= 1'b1;
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	fval �½��ؼĴ���
	//	1.�������ؼĴ�����Чʱ����fval�½��ص�ʱ�򣬼Ĵ�����1
	//	2.�������ؼĴ�����Чʱ���Ĵ�������
	//	3.�������أ����½��ص�˳��
	//	4.�������غ��½��ؼĴ�������Ч��ʱ��˵����ʹ����Ч��ʱ�򣬾���һ������֡
	//	5.��������ɿ���֮�󣬵�һ֡��3aͳ�Ʋ������жϡ�Ŀ����Ϊ�˷�ֹ���ɺ�ĵ�һ֡���ܻ��ǲ�֡������ͳ�ƴ���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(fval_rise_reg) begin
			if(fval_fall) begin
				full_frame_state	<= 1'b1;
			end
		end
		else begin
			full_frame_state	<= 1'b0;
		end
	end

	//  ===============================================================================================
	//	ref ***�ڲ��ж�״̬***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	--ref 2a-�ڲ��ж�״̬
	//	1.����֡ʹ����Чʱ���ڲ��ж�״̬��������
	//	2.����֡ʹ����Чʱ���ж�ʹ����Ч���ڲ��ж�״̬����
	//	3.����֡ʹ����Чʱ���ж�ʹ����Ч���ڳ��ź��½���(��һ��֮����ź�)ʱ���ڲ��ж�״̬��1
	//	4.����֡ʹ����Чʱ���ж�ʹ����Ч��clear��Чʱ���ڲ��ж�״̬����
	//	5.3 4 ͬʱ������3����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!full_frame_state) begin
			internal_state[0]	<= 1'b0;
		end
		else begin
			if(!i_interrupt_en_grey) begin
				internal_state[0]	<= 1'b0;
			end
			else begin
				if(fval_fall_dly0) begin
					internal_state[0]	<= 1'b1;
				end
				else if(iv_interrupt_clear[0]) begin
					internal_state[0]	<= 1'b0;
				end
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	--ref wb-�ڲ��ж�״̬
	//	1.����֡ʹ����Чʱ���ڲ��ж�״̬��������
	//	2.����֡ʹ����Чʱ���ж�ʹ����Ч���ڲ��ж�״̬����
	//	3.����֡ʹ����Чʱ���ж�ʹ����Ч���ڳ��ź��½���(��һ��֮����ź�)ʱ���ڲ��ж�״̬��1
	//	4.����֡ʹ����Чʱ���ж�ʹ����Ч��clear��Чʱ���ڲ��ж�״̬����
	//	5.3 4 ͬʱ������3����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!full_frame_state) begin
			internal_state[1]	<= 1'b0;
		end
		else begin
			if(!i_interrupt_en_wb) begin
				internal_state[1]	<= 1'b0;
			end
			else begin
				if(fval_fall_dly0) begin
					internal_state[1]	<= 1'b1;
				end
				else if(iv_interrupt_clear[1]) begin
					internal_state[1]	<= 1'b0;
				end
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	ref ***�ӿ��ж�״̬***
	//	1.�ڲ��ж�״̬����ʱ���ӿ��ж�״̬����
	//	2.�ڲ��ж�״̬=1ʱ����int������ʱ���ӿ��ж�״̬=1
	//  -------------------------------------------------------------------------------------
	genvar j;
	generate
		for(j=0;j<=1;j=j+1) begin
			always @ (posedge clk) begin
				if(!internal_state[j]) begin
					interface_state[j]	<= 1'b0;
				end
				else begin
					if(int_rise) begin
						interface_state[j]	<= 1'b1;
					end
				end
			end
		end
	endgenerate
	assign	ov_interrupt_state	= interface_state;

	//  ===============================================================================================
	//	ref ***50ms �жϼ��**
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	-- ref 50ms������
	//	1.72MHz��ʱ�ӣ���Ҫ������3600000���Ż���50ms��16������0x36EE80��22λ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(int_rise) begin
			div_time_interval_cnt	<= 'b0;
		end
		else begin
			if(div_time_interval_cnt==TIME_INTERVAL) begin
				div_time_interval_cnt	<= div_time_interval_cnt;
			end
			else begin
				div_time_interval_cnt	<= div_time_interval_cnt + 1'b1;
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	����ʱ�䵽��־
	//	1.����������50msʱ��time up=1
	//	2.������δ����50msʱ��time up=0
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(div_time_interval_cnt==TIME_INTERVAL) begin
			time_up	<= 1'b1;
		end
		else begin
			time_up	<= 1'b0;
		end
	end

	//  -------------------------------------------------------------------------------------
	//	--ref �жϷ�����־
	//	1.��50msʱ�䵽�ˣ���fval�½���(������֮����ź�)��Ч������ж�״̬ʱȫ�㣬�����Ϊ0
	//	2.��50msʱ�䵽�ˣ���fval�½���(������֮����ź�)��Ч������ж�״̬ʱ������1��1�������Ϊ1
	//	3.�����жϱ�־=0
	//	4.�жϱ�־�ߵ�ƽ�����1��ʱ������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(time_up&fval_fall_dly1) begin
			if(internal_state[1:0]==2'b00) begin
				int_rise	<= 1'b0;
			end
			else begin
				int_rise	<= 1'b1;
			end
		end
		else begin
			int_rise	<= 1'b0;
		end
	end

	//  ===============================================================================================
	//	ref ***�����ж�***
	//	3014���ж��ź��Ǹ���Ч����Ϳ����100ns
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	�ж�չ��Ĵ���
	//	1.���жϱ�־��Чʱ��չ��Ĵ�������
	//	2.���жϱ�־��Чʱ��������������λ=1����ֹͣ�����������������
	//	3.72MHz��Ƶ�ʣ�����16�����ڣ������222ns
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(int_rise) begin
			extend_int_cnt	<= 5'b0;
		end
		else begin
			if(extend_int_cnt[4]==1'b1) begin
				extend_int_cnt	<= extend_int_cnt;
			end
			else begin
				extend_int_cnt	<= extend_int_cnt + 1'b1;
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	�жϼĴ�������չ��Ĵ������λȡ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		interrupt_reg	<= !extend_int_cnt[4];
	end
	assign	o_interrupt	= interrupt_reg;



endmodule