//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : strobe_filter
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/1/12 17:13:14	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ��strobe�ź��˲���MT9P031���ع��ź���bug����Ҫ�����˲�
//              1)  : ��strobe���С�ڵ���1�п��ʱ�����ܷ���strobe�ź�
//
//              2)  : ��strobe��ȴ���1�п��ʱ���������strobe�ź�
//
//              3)  : �����strobe�źſ�Ȳ��䣬λ�����Ų��1��
//
//              4)  : ��ģ���ڲ�ͳ���п�ȣ�����lval���첽ʱ�����п����ٲ���1������Ҫע��˴�
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module strobe_filter (
	input				clk						,	//����ʱ�ӣ�72MHz
	input				i_acquisition_start		,	//�����źţ�0-ͣ�ɣ�1-����
	input				i_stream_enable			,	//��ʹ���źţ�0-ͣ�ɣ�1-����
	input				i_fval					,	//����Ч�źţ��첽�źţ���i_lval���ض���
	input				i_lval					,	//����Ч�źţ��첽�źţ���i_fval���ض���
	input				i_sensor_strobe			,	//�ع��źţ��첽�źţ����ع��źſ��С��1��ʱ����������ع��ź�
	output	[12:0]		ov_strobe_length_reg	,	//������strobe���
	output				o_strobe_filter				//�����˲�����ع��ź�
	);

	//	ref signals
	reg		[1:0]		fval_shift				= 2'b0;
	reg		[3:0]		lval_shift				= 4'b0;
	wire				lval_rise				;
	reg		[1:0]		strobe_shift			= 2'b0;
	wire				strobe_int				;
	reg		[1:0]		lval_rise_cnt			= 2'b0;
	wire				lperiod_length_upload	;
	reg		[12:0]		lperiod_length_cnt		= 13'h0000;
	reg		[12:0]		lperiod_length_reg		= 13'h1fff;
	reg		[12:0]		strobe_length_reg		= 13'h1fff;
	reg		[12:0]		strobe_length_cnt		= 13'h0000;
	reg					enable					= 1'b0;
	reg					strobe_dout				= 1'b0;



	//	ref ARCHITECTURE
	//  ===============================================================================================
	//	ref �첽�źſ�ʱ������
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	fval ������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_shift	<= {fval_shift[0],i_fval};
	end

	//  -------------------------------------------------------------------------------------
	//	lval �����ģ���Ϊfval��lval�Ǳ��ض���ģ�Ҫ��fval=1��ʱ����lval�������أ���Ҫ��lva����ʱ2��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		lval_shift	<= {lval_shift[2:0],i_lval};
	end
	assign	lval_rise	= (lval_shift[3]==1'b0 && lval_shift[2]==1'b1) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//	strobe ������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		strobe_shift	<= {strobe_shift[0],i_sensor_strobe};
	end

	//	-------------------------------------------------------------------------------------
	//	���strobe�źų�����fval=1֮�ڣ���Ҫ�˵��ġ�
	//	1.�Ӳ��Խ���������strobe������fval=1֮�ڣ��϶���1�еĿ�ȡ�
	//	2.�������ε�Ŀ������ǿ�˲��Ľ�׳��
	//	-------------------------------------------------------------------------------------
	assign	strobe_int	= (fval_shift[1]==1'b1) ? 1'b0 : strobe_shift[1];

	//  ===============================================================================================
	//	ref �����ڼ�������fval=1��ʱ�����
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	lval�����ظ���������
	//	1.��fval=0ʱ,����������
	//	2.����fval=1��lval�����ص���ʱ,cnt++
	//	3.��lval cnt����������1'b1ʱ,����������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!fval_shift[1]) begin
			lval_rise_cnt	<= 2'b0;
		end
		else begin
			if(lval_rise) begin
				if(lval_rise_cnt==2'b10) begin
					lval_rise_cnt	<= lval_rise_cnt;
				end
				else begin
					lval_rise_cnt	<= lval_rise_cnt + 1'b1;
				end
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	��lval rise cnt��lval rise������1ʱ��upload��־=1.
	//	1.��ʱ˵����fval=1�ڼ��Ѿ�����2��lval��������
	//  -------------------------------------------------------------------------------------
	assign	lperiod_length_upload	= (lval_rise_cnt==2'b01 && lval_rise==1'b1) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//	�����ڼ�����
	//	1.��lval rise cnt=0ʱ�������ڼ���������
	//	2.��lval rise cnt=1ʱ�������ڼ�����++
	//	3.��lval rise cnt=1ʱ����������ڼ�����ȫ1,����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(lval_rise_cnt==2'b0) begin
			lperiod_length_cnt	<= 'b0;
		end
		else if(lval_rise_cnt==2'b01) begin
			if(lperiod_length_cnt==13'h1ff0) begin
				lperiod_length_cnt	<= lperiod_length_cnt;
			end
			else begin
				lperiod_length_cnt	<= lperiod_length_cnt + 1'b1;
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	�����ڼĴ���
	//	1.�������ź���Чʱ�������µ������ڳ����Ѿ�����������Ĵ���=������+15���˴���10��Ϊ�˱�֤1�п�ȵ�strobeҲ�ᱻ�˵�
	//	2.�����ڼĴ����ϵ��ʼֵ��ȫ1��Ϊ����Sensor��һ֡�����fval=1��ʼʱ����strobe����������󴥷������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(lperiod_length_upload) begin
			lperiod_length_reg	<= lperiod_length_cnt+4'hf;
		end
	end
	
	//  ===============================================================================================
	//	ref strobe �˲�
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	strobe �˲����ȼĴ���
	//	1.��strobe ���ȼ���������ʱ�����ܸ��� strobe ���ȼĴ���
	//	2.strobe���ȼĴ����ϵ��ʼֵ��ȫ1��Ϊ����Sensor��һ֡�����fval=1��ʼʱ����strobe����������󴥷������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(strobe_length_cnt==13'h0000) begin
			strobe_length_reg	<= lperiod_length_reg;
		end
	end
	assign	ov_strobe_length_reg	= strobe_length_reg;
	
	//  -------------------------------------------------------------------------------------
	//	strobe �˲����ȼ�����
	//	1.��strobe�����0ʱ�����strobe������1���������++�����������=�Ĵ������򱣳�
	//	2.��strobe�����0ʱ�����strobe������0�������������
	//	3.��strobe�����1ʱ�����strobe������1�������������
	//	4.��strobe�����1ʱ�����strobe������0���������--�����������=ȫ0���򱣳�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!strobe_dout) begin
			if(strobe_int) begin
				if(strobe_length_cnt==strobe_length_reg) begin
					strobe_length_cnt	<= strobe_length_cnt;
				end
				else begin
					strobe_length_cnt	<= strobe_length_cnt + 1'b1;
				end
			end
			else begin
				strobe_length_cnt	<= 13'b0;
			end
		end
		else begin
			if(strobe_int) begin
				strobe_length_cnt	<= strobe_length_cnt;
			end
			else begin
				if(strobe_length_cnt==13'h0000) begin
					strobe_length_cnt	<= strobe_length_cnt;
				end
				else begin
					strobe_length_cnt	<= strobe_length_cnt - 1'b1;
				end
			end
		end
	end

	//  ===============================================================================================
	//	ref ���
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	ʹ���ź�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		enable	<= i_stream_enable&i_acquisition_start;
	end

	//  -------------------------------------------------------------------------------------
	//	strobe���
	//	1.���ʹ����Ч���������Ϊ0
	//	2.���ʹ����Ч����strobe������1�����˲��������ﵽ���˲��Ĵ����ĳ��ȣ����1
	//	3.���ʹ����Ч����strobe������0�����˲��Ĵ���=ȫ�㣬���0
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!enable) begin
			strobe_dout	<= 1'b0;
		end
		else begin
			if(strobe_int==1'b1 && strobe_length_cnt==strobe_length_reg) begin
				strobe_dout	<= 1'b1;
			end
			else if(strobe_int==1'b0 && strobe_length_cnt==13'h0000) begin
				strobe_dout	<= 1'b0;
			end
		end
	end

	assign	o_strobe_filter	= strobe_dout;


endmodule
