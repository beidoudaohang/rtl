//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : testcase_1
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/4/10 16:50:28	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ���ڴ�С��16x16�������ź���Ч������ģʽ�µ�����״��
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`include 	"SHARP_RJ33B4_DEF.v"
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module testcase_1 ();

	//	ref signals
	//	===============================================================================================
	//	--ref parameter
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	TESTCASE
	//	-------------------------------------------------------------------------------------
	parameter	TESTCASE_NUM			= "testcase_1"			;	//����ģ����Ҫʹ���ַ���
	//	-------------------------------------------------------------------------------------
	//	sensor model parameter
	//	-------------------------------------------------------------------------------------


	//	-------------------------------------------------------------------------------------
	//	dut paramter
	//	-------------------------------------------------------------------------------------


	//	-------------------------------------------------------------------------------------
	//	monitor paramter
	//	-------------------------------------------------------------------------------------

	//	-------------------------------------------------------------------------------------
	//	testcase parameter
	//	-------------------------------------------------------------------------------------
//	parameter	CLK_PERIOD				= 22.222	;	//ʱ��Ƶ�ʣ�45MHz
	parameter	CLK_PERIOD				= 16.667	;	//ʱ��Ƶ�ʣ�60MHz
//	parameter	CLK_PERIOD				= 20.833	;	//ʱ��Ƶ�ʣ�48MHz

	//	===============================================================================================
	//	--ref signal
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	sensor signal
	//	-------------------------------------------------------------------------------------

	//	-------------------------------------------------------------------------------------
	//	dut signal
	//	-------------------------------------------------------------------------------------
	reg								clk					= 1'b0	;
	reg								reset				= 1'b0	;
	reg								i_start_acquisit	= 1'b1	;
	reg								i_trigger			= 1'b0	;
	reg								i_triggermode		= 1'b0	;
	reg		[`LINE_WD - 1:0]		iv_href_start		= 'b0	;
	reg		[`LINE_WD - 1:0]		iv_href_end			= 'b0	;
	reg		[`LINE_WD - 1:0]		iv_hd_rising		= 'b0	;
	reg		[`LINE_WD - 1:0]		iv_hd_falling		= 'b0	;
	reg		[`LINE_WD - 1:0]		iv_sub_rising		= 'b0	;
	reg		[`LINE_WD - 1:0]		iv_sub_falling		= 'b0	;
	reg		[`FRAME_WD - 1:0]		iv_vd_rising		= 'b0	;
	reg		[`FRAME_WD - 1:0]		iv_vd_falling		= 'b0	;
	reg		[`EXP_WD - 1:0]			iv_xsg_width		= 'b0	;

	reg								i_ad_parm_valid		= 1'b0	;

	//	ref ARCHITECTURE

	//	===============================================================================================
	//	ref ***tb ��ģ�鼤��***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	--ref Sensor
	//	-------------------------------------------------------------------------------------
	always	#(CLK_PERIOD/2.0)	clk	= !clk;

	//	-------------------------------------------------------------------------------------
	//	--ref DUT
	//	-------------------------------------------------------------------------------------

	//	-------------------------------------------------------------------------------------
	//	--ref ����ʱ��
	//	-------------------------------------------------------------------------------------
	initial begin
		#200
		//		repeat(20) @ (negedge harness.o_fval);
		//		repeat(30) @ (negedge driver_mt9p031.o_fval);
		#20000
		#40000000
		$stop;
	end

	//	===============================================================================================
	//	ref ***����bfm task***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	��λ
	//	-------------------------------------------------------------------------------------
	initial begin
		reset 			= 1;
		#200 reset 		= 0;
	end

	//	-------------------------------------------------------------------------------------
	//	����ccd����
	//	-------------------------------------------------------------------------------------
	//	-------------------------------------------------------------------------------------
	//	�̶�λ��
	//	-------------------------------------------------------------------------------------
	initial begin
		iv_hd_rising			= `HD_RISING	;
		iv_hd_falling			= `HD_FALLING	;
		iv_vd_rising			= `VD_RISING	;
		iv_vd_falling			= `VD_FALLING	;
		iv_sub_rising			= `SUB_RISING	;
		iv_sub_falling			= `SUB_FALLING	;
	end

	initial begin
		iv_href_start			= `HREF_START_DEFVALUE		;
		iv_href_end				= `HREF_END_DEFVALUE		;
	end

	//	-------------------------------------------------------------------------------------
	//	����ccd�ع�ʱ��
	//	-------------------------------------------------------------------------------------
	initial begin
		iv_xsg_width			= `XSG_WIDTH	;
	end


	initial begin
//		harness.bfm_ccd.readout_reg_cfg(0,0,1292,964);
		harness.bfm_ccd.readout_reg_cfg(0,0,660,492);
//		harness.bfm_ccd.readout_reg_cfg(8,960);
//		harness.bfm_ccd.exp_time_us(40);
//		harness.bfm_ccd.exp_time_us(50);
//		harness.bfm_ccd.exp_time_us(100);
//		harness.bfm_ccd.exp_time_us(20);
//		harness.bfm_ccd.exp_time_us(41076);
//		harness.bfm_ccd.exp_time_us(49736);
		harness.bfm_ccd.exp_time_us(1000);
	end


	initial begin
		i_start_acquisit		= 1'b0	;
		#10000
		i_start_acquisit		= 1'b1	;
	end



endmodule
