//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : led_ctrl
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/12/1 14:54:14	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : led ����ƿ���ģ��
//              1)  : ���ݼĴ�����������������ⲿ��LED��״̬
//
//              2)  : �ⲿ��2��LED����ƺ��̵ƣ��ߵ�ƽ�����������ƶ���ʱ��Ϊ��ɫ
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module led_ctrl # (
	parameter		LED_CTRL_WIDTH					= 5		//LED CTRL �Ĵ������
	)
	(
	//ʱ��
	input								clk				,	//ʱ���ź�
	//�Ĵ����ź�
	input								i_usb_slwr_n	,	//GPIF д�źţ�clk_gpifʱ����
	//  -------------------------------------------------------------------------------------
	//	led_ctrl
	//	0x00:��Ƴ�������ʱFPGA����δ��ɼ��ػ����������С�
	//	0x01:�����ݴ���ʱ���̵Ƴ�������ͼ�����ݴ���ʱ���̵���˸����ͼ������ʱϨ����ͼ������ʱ������
	//	0x10:�Ƶ���˸(1Hz)����ʱ������һ����󣬱����û���������ʧ�ܡ�
	//  -------------------------------------------------------------------------------------
	input	[LED_CTRL_WIDTH-1:0]		iv_led_ctrl		,	//led���ƼĴ�����FPGA�ⲿ���Ӻ�������LED�ƣ�����LEDͬʱ��ʱΪ��ɫ��
	//FPGA ����
	output								o_f_led_gre		,	//��ɫָʾ�ƣ��ߵ�ƽ����
	output								o_f_led_red			//��ɫָʾ�ƣ��ߵ�ƽ����
	);

	//	ref signals
	reg		[1:0]		usb_wr_shift	= 2'b0;
	reg		[4:0]		led_ctrl_reg	= 5'b0;
	reg		[25:0]		div_72m_1hz_cnt	= 26'b0;
	reg					twinkle_1hz		= 1'b0;
	reg					led_gre			= 1'b0;
	reg					led_red			= 1'b0;

	//	-------------------------------------------------------------------------------------
	//	����׶Σ�LED��˸������50ms
	//	-------------------------------------------------------------------------------------
	reg		[21:0]		transit_twinkle_period		= 22'h35ee80;
	reg					twinkle_20hz_cnt_en			= 1'b0;
	reg		[21:0]		div_72m_20hz_cnt			= 22'b0;
	reg					twinkle_20hz				= 1'b0;


	//	ref ARCHITECTURE
	//	===============================================================================================
	//	ref ***led_ctrl***
	//	===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	��ʱ����ͬ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		usb_wr_shift	<= {usb_wr_shift[0],i_usb_slwr_n};
	end

	//	-------------------------------------------------------------------------------------
	//	����led_ctrl�Ĵ���
	//	����Ϊ�Ƿ�ֵʱ��led_ctrl_reg���ܸ���
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		case(iv_led_ctrl[4:0])
			5'h00,5'h01,5'h10	: begin
				led_ctrl_reg	<= iv_led_ctrl;
			end
			default	: begin
				led_ctrl_reg	<= led_ctrl_reg;
			end
		endcase
	end

	//  -------------------------------------------------------------------------------------
	//	1Hz�ź�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(div_72m_1hz_cnt==26'h22550FF) begin
			div_72m_1hz_cnt	<= 26'b0;
		end
		else begin
			div_72m_1hz_cnt	<= div_72m_1hz_cnt + 1'b1;
		end
	end

	always @ (posedge clk) begin
		if(div_72m_1hz_cnt==26'h22550FF) begin
			twinkle_1hz	<= !twinkle_1hz;
		end
	end

	//  -------------------------------------------------------------------------------------
	//	�̵�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		case(led_ctrl_reg[4:0])
			5'h00 	: led_gre	<= 1'b0;
			5'h01	: led_gre	<= twinkle_20hz;
			5'h10	: led_gre	<= twinkle_1hz;
			default	: ;//��Ҫ���û����ȷ˵����������Ŀǰ��ȡ����ǵĴ�����
		endcase
	end
	assign	o_f_led_gre	= led_gre;

	//  -------------------------------------------------------------------------------------
	//	���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		case(led_ctrl_reg[4:0])
			5'h00	: led_red	<= 1'b1;
			5'h01	: led_red	<= 1'b0;
			5'h10	: led_red	<= twinkle_1hz;
			default	: ;//��Ҫ���û����ȷ˵����������Ŀǰ��ȡ����ǵĴ�����
		endcase
	end
	assign	o_f_led_red	= led_red;

	//	===============================================================================================
	//	ref ***����׶���˸***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	������ʹ��
	//	1.������50msʱ���ӷ���ʹ��ȡ��
	//	2.��������û�м�����50msʱ��ֻҪд�ź���Ч��������ʹ�ܾ���Ч
	//	3.һ��д�ź���Ч��������ʹ�ܾ���Ч��һ���������ӵ����ֵ��������ʹ��ȡ��
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(div_72m_20hz_cnt==transit_twinkle_period) begin
			twinkle_20hz_cnt_en	<= 1'b0;
		end
		else if(!usb_wr_shift[1]) begin
			twinkle_20hz_cnt_en	<= 1'b1;
		end
	end

	//	-------------------------------------------------------------------------------------
	//	div_72m_20hz_cnt ��˸������
	//	1.���������ӵ�50ms������0
	//	2.�ڼ�����û�е������ֵʱ��ֻҪ������ʹ����Ч��������
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(div_72m_20hz_cnt==transit_twinkle_period) begin
			div_72m_20hz_cnt	<= 22'b0;
		end
		else if(twinkle_20hz_cnt_en) begin
			div_72m_20hz_cnt	<= div_72m_20hz_cnt + 1'b1;
		end
	end

	//	-------------------------------------------------------------------------------------
	//	��˸�ź�
	//	1.����������0ʱ����˸�ź�Ϊ1��������led
	//	2.�����������ӵ�1/4����ʱ��Ϩ��led
	//	3.�ߵ�ƽʱ��ֻ��1/4���ڣ�led����ʱ��϶�
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(div_72m_20hz_cnt==22'b0) begin
			twinkle_20hz	<= 1'b1;
		end
		else if(div_72m_20hz_cnt=={2'b00,transit_twinkle_period[21:2]}) begin
			twinkle_20hz	<= 1'b0;
		end
	end


endmodule
