//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : bfm
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/4/8 11:28:42	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------
module bfm # (
	parameter		DATA_WIDTH			= 32		,	//���ݿ��
	parameter		PTR_WIDTH			= 2			,	//��дָ���λ��1-���2֡ 2-���4֡ 3-���8֡ 4-���16֡ 5-���32֡
	parameter		FRAME_SIZE_WIDTH	= 25			//һ֡��Сλ����DDR3��1Gbitʱ�����������128Mbyte����mcb p3 ��λ����32ʱ��25λ���size���������㹻��
	)
	();

	//	ref signals
	//	-------------------------------------------------------------------------------------
	//	�����ź�
	//	-------------------------------------------------------------------------------------
	reg		[PTR_WIDTH-1:0]				iv_frame_depth			;
	reg									i_start_full_frame		= 1'b1;
	reg									i_start_quick			= 1'b1;
	wire	[FRAME_SIZE_WIDTH-1:0]		iv_frame_size			;
	reg		[31:0]						iv_transfer_count		= 32'b0;
	reg		[31:0]						iv_transfer_size		= 32'b0;
	reg		[31:0]						iv_transfer1_size		= 32'b0;
	reg		[31:0]						iv_transfer2_size		= 32'b0;



	//	ref ARCHITECTURE

	//  ===============================================================================================
	//	ref ***֡�� task***
	//  ===============================================================================================
	task frame_depth;
		input	[PTR_WIDTH-1:0]		iv_frame_depth_input;
		begin
			#1
			iv_frame_depth	= iv_frame_depth_input;
		end
	endtask

	//	-------------------------------------------------------------------------------------
	//	֡���С
	//	-------------------------------------------------------------------------------------
	assign	iv_frame_size		= (driver_mt9p031.bfm_mt9p031.iv_line_active_pix_num * driver_mt9p031.bfm_mt9p031.iv_line_active_num);

	//	-------------------------------------------------------------------------------------
	//	start_ff
	//	-------------------------------------------------------------------------------------
	task start_ff_high;
		begin
			#1
			i_start_full_frame	= 1'b1;
		end
	endtask
	
	task start_ff_low;
		begin
			#1
			i_start_full_frame	= 1'b1;
		end
	endtask

	//	-------------------------------------------------------------------------------------
	//	start_qk
	//	-------------------------------------------------------------------------------------
	task start_qk_high;
		begin
			#1
			i_start_quick	= 1'b1;
		end
	endtask
	
	task start_qk_low;
		begin
			#1
			i_start_quick	= 1'b1;
		end
	endtask

	//	-------------------------------------------------------------------------------------
	//	si info
	//	-------------------------------------------------------------------------------------
	task si_info;
		begin
			#1
			iv_transfer_size	= 32'h100000;
			#1
			iv_transfer_count	= iv_frame_size/iv_transfer_size;
			#1
			iv_transfer1_size	= (((iv_frame_size-iv_transfer_size*iv_transfer_count)/32'h400)*32'h400);
			#1
			if((iv_frame_size-iv_transfer_size*iv_transfer_count-iv_transfer1_size)!=0) begin
				iv_transfer2_size	= 32'h400;
			end
			else begin
				iv_transfer2_size	= 32'h0;
			end
		end
	endtask




endmodule
