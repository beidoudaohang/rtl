//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : trigger_extend
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/12/2 17:20:57	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :չ��ģ�飬����Sensor�Ĵ����źŶԵ͵�ƽʱ����Ҫ��trigger����Ҫ1�е�ʱ���ȣ�8192�������
//              1)  : �����ź���1��ʱ�ӿ�ȵĸ�����
//
//              2)  : ����ź���չ��Ϊ8192��ȵĵ�����
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module trigger_extend (
	input			clk					,	//ʱ��
	//�Ĵ���
	input			i_trigger_mode		,	//����ģʽ��0-����ģʽ��1-����ģʽ
	input			i_stream_enable		,	//��ʹ���ź�
	input			i_acquisition_start	,	//�����źţ�0-ͣ�ɣ�1-����
	//�����ź�
	input			i_din				,	//���봥���ź�
	output			o_dout_n				//��������źţ��͵�ƽ��Ч
	);

	//	ref signals
	parameter				EXTEND_LENGTH	= 8192;	//Ҫչ��ĳ���
	reg						enable			= 1'b0;
	reg						extending		= 1'b0;
	reg		[12:0]			extend_cnt		= 13'b0;
	reg						dout_reg		= 1'b1;
	

	//	ref ARCHITECTURE

	//  -------------------------------------------------------------------------------------
	//	ʹ���źţ���ioͨ�������1��ģ�����������
	//	1.������ʹ���źŶ�ʹ��ʱ�����1
	//	2.������ʹ���ź���1����0ʱ�����0
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		enable	<= i_trigger_mode&i_stream_enable&i_acquisition_start;
	end

	//  -------------------------------------------------------------------------------------
	//	����չ��ı�־
	//	1.��չ���������չ�������ʱ�����0
	//	2.�������ź���1��ʹ����Чʱ�����1����ʼչ��
	//	3.ʹ���źŲ�����������չ����ź�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(extend_cnt==EXTEND_LENGTH-1) begin
			extending	<= 1'b0;
		end
		else if(i_din==1'b1 && enable==1'b1) begin
			extending	<= 1'b1;
		end
	end

	//  -------------------------------------------------------------------------------------
	//	չ�������
	//	1.��չ���������չ�������ʱ��չ�����������
	//	2.������չ���־=1ʱ��չ�������+1
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(extend_cnt==EXTEND_LENGTH-1) begin
			extend_cnt	<= 13'b0;
		end
		else if(extending) begin
			extend_cnt	<= extend_cnt + 1'b1;
		end
	end

	//  -------------------------------------------------------------------------------------
	//	���ȡ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		dout_reg	<= !extending;
	end
	assign	o_dout_n	= dout_reg;


endmodule
