//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : trailer
//  -- �����       : ��ǿ
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- ��ǿ         :| 2014/12/3 16:50:10	:|  ���ݼ���Ԥ������
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������
//              1)  : U3V��ʽtrailerģ�飬��ϳɷ���U3V��ʽtrailer��
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module trailer # (
	parameter				DATA_WD						= 32	,	//�����������λ������ʹ��ͬһ���
	parameter				SHORT_REG_WD 				= 16	,	//�̼Ĵ���λ��
	parameter				REG_WD 						= 32	,	//�Ĵ���λ��
	parameter				LONG_REG_WD 				= 64		//���Ĵ���λ��
	)
	(
//  ===============================================================================================
//  ��һ���֣�ʱ�Ӹ�λ
//  ===============================================================================================
	input							reset						,	//��λ�źţ��ߵ�ƽ��Ч������ʱ��ʱ����
	input							clk							,	//ʱ���źţ�����ʱ��ʱ����ͬ�ڲ�����ʱ��
//  ===============================================================================================
//  �ڶ����֣�β����־
//  ===============================================================================================
	input							i_trailer_flag				,	//ͷ����־
//  ===============================================================================================
//  �������֣����ƼĴ�����chunk��Ϣ��ֻ���Ĵ���
//  ===============================================================================================
	input							i_chunk_mode_active			,	//chunk�ܿ��أ����ش�Payload Typeʹ��Ϊimage extend chunk ���ͣ�chunk�ر�Ϊimage����
	input							i_chunkid_en_ts	    		,	//ʱ���chunkʹ��
    input							i_chunkid_en_fid	        ,   //frame id chunkʹ��
	input		[LONG_REG_WD-1  :0]	iv_blockid					,	//ͷ����chunk��β����blockid��Ϣ����һ֡��block ID��0��ʼ��������һ֡block IDΪ0
	input		[SHORT_REG_WD-1 :0]	iv_status					, 	//β���еĵ�ǰ֡״̬
	input		[REG_WD-1		:0]	iv_valid_payload_size		, 	//β���е���Ч���ش�С�ֶ�
	input		[SHORT_REG_WD-1 :0]	iv_trailer_size_y			, 	//β���е���Ч�߶��ֶ�
//  ===============================================================================================
//  ���Ĳ��֣��С�������Ч������
//  ===============================================================================================
	output	reg						o_data_valid				,	//�����ͷβ��������Ч�ź�
	output	reg	[DATA_WD-1:0]		ov_data							//
	);

//  ===============================================================================================
//  ���ز���
//  ===============================================================================================
	localparam						TRAILER_LENTH	=	4'd9	;	//β������9
//  ===============================================================================================
//  �����ͼĴ�������
//  ===============================================================================================
	reg			[3				:0]	count          = 	4'h0	;	//���������������β���е��ź�
	reg								chunk_mode_active_r			;	//
	reg								chunkid_en_ts_r	            ;	//
	reg								chunkid_en_fid_r            ;	//
	reg			[7				:0]	chunk_layout_id	=	8'h0 	;
//  ===============================================================================================
//  chunk_layoutid�仯
//  ===============================================================================================
	always @ (posedge clk)
		begin
			chunk_mode_active_r	<=   i_chunk_mode_active	;
			chunkid_en_ts_r	    <=   i_chunkid_en_ts		;
			chunkid_en_fid_r    <=   i_chunkid_en_fid	    ;
		end

	always @ (posedge clk)
		begin
			if ( (chunk_mode_active_r ^ i_chunk_mode_active) || (chunkid_en_ts_r ^ i_chunkid_en_ts) || (chunkid_en_fid_r ^ i_chunkid_en_fid))
				chunk_layout_id	<= chunk_layout_id +1;
		end
//  ===============================================================================================
//  i_trailer_flag�ڼ���
//  ===============================================================================================
	always @ (posedge clk) begin
		if(i_trailer_flag) begin
			count	<=	count + 4'h1;
		end
		else begin
			count	<=	4'h0;
		end
	end
//  -------------------------------------------------------------------------------------
//  ����trailer�����ݣ�����ʽ����Image Extended Chunk Trailer��ʽ
//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if ( reset ) begin
			ov_data <= 	32'h0;
		end
		else begin
			case ( count )
				4'h1	:	ov_data	<=	32'h54563355				;
				4'h2	:   ov_data	<=	{13'h4,i_chunk_mode_active,2'b00,16'd0}	;	//����ʹ��λ����һ��ƴ�ӣ���i_chunk_mode_activeʹ�ܣ�����Ϊ36������Ϊ32
				4'h3	:   ov_data	<=	iv_blockid[31:0]          	;
				4'h4	:   ov_data	<=	iv_blockid[63:32]         	;
				4'h5	:   ov_data	<=	{16'h00,iv_status}			;				//����ֻ֧��Image��0x0001����Image Extended Chunk��0x4001��
				4'h6	:   ov_data	<=	iv_valid_payload_size[31:0]	;
				4'h7	:   ov_data	<=	32'h0						;
				4'h8	:   ov_data	<=	{16'h00,iv_trailer_size_y}	;
				4'h9	:   ov_data	<=	{24'h0,chunk_layout_id}		;				//chunk_layout_idΪ0
				default	:  	ov_data <= 	32'h0						;
			endcase
		end
	end
//  -------------------------------------------------------------------------------------
//  ���o_data_valid�ź�,i_chunk_mode_active��Чʱ9��ʱ�ӿ�ȣ���Чʱ8��ʱ�ӿ��
//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if ( reset ) begin
			o_data_valid	<=	1'b0;
		end
		else if ( count == 4'h1 )begin
			o_data_valid	<=	1'b1;
		end
		else if ( (count == TRAILER_LENTH) && (~i_chunk_mode_active)  ) begin
			o_data_valid	<=	1'b0;
		end
		else if ( (count == TRAILER_LENTH+1) && i_chunk_mode_active  ) begin
			o_data_valid	<=	1'b0;
		end
	end

endmodule