//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : gen_wr_data
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/6/9 16:25:06	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//`include			"gen_wr_data_def.v"
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module gen_wr_data (
	input			clk		,
	//	input			reset	,
	output	[31:0]	ov_image_data

	);

	//	ref signals

	reg		[7:0]	lfsr 	= 8'hab;

	//	ref ARCHITECTURE


	always @ (posedge clk) begin
		lfsr[0]	<= lfsr[7];
		lfsr[1]	<= lfsr[6];
		lfsr[2]	<= lfsr[5]^lfsr[4];
		lfsr[3]	<= lfsr[4]^lfsr[3];
		lfsr[4]	<= lfsr[3]^lfsr[2];
		lfsr[5]	<= lfsr[2]^lfsr[1];
		lfsr[6]	<= lfsr[1];
		lfsr[7]	<= lfsr[0];
	end

	assign	ov_image_data	= {4{lfsr}};

endmodule
