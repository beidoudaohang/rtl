//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : cs_top
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/6/5 14:45:18	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//`include			"cs_top_def.v"
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module cs_top (
	input			CLK			,
	input	[119:0]	TRIG0		,
	input	[31:0]	ASYNC_IN	,
	output	[31:0]	ASYNC_OUT
	);

	//	ref signals

	wire	[35:0]	CONTROL0;
	wire	[35:0]	CONTROL1;

	//	ref ARCHITECTURE

	chipscope_icon chipscope_icon_inst (
	.CONTROL0	(CONTROL0	),
	.CONTROL1	(CONTROL1	)
	);

	chipscope_ila chipscope_ila_inst (
	.CONTROL	(CONTROL0	),
	.CLK		(CLK		),
	.TRIG0		(TRIG0		)
	);

	chipscope_vio chipscope_vio_inst (
	.CONTROL	(CONTROL1	),
	.ASYNC_IN	(ASYNC_IN	),
	.ASYNC_OUT	(ASYNC_OUT	)
	);




endmodule
