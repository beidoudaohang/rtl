//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : testcase_14
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/4/10 16:50:28	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : fval��С���� ��С��3
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module testcase_14 ();

	//	ref signals
	//	===============================================================================================
	//	--ref parameter
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	TESTCASE
	//	-------------------------------------------------------------------------------------
	parameter	TESTCASE_NUM			= "testcase_14"			;	//����ģ����Ҫʹ���ַ���
	//	-------------------------------------------------------------------------------------
	//	sensor model parameter
	//	-------------------------------------------------------------------------------------
	parameter	IMAGE_SRC				= "RANDOM"				;	//"RANDOM" or "FILE" or "LINE_INC" or "FRAME_INC"
	parameter	DATA_WIDTH				= 10					;	//8 10 12 max is 16
	parameter	CHANNEL_NUM				= 4						;	//ͨ����
	parameter	SENSOR_CLK_DELAY_VALUE	= 3						;	//Sensor оƬ�ڲ���ʱ ��λns
	parameter	CLK_DATA_ALIGN			= "RISING"				;	//"RISING" - ���ʱ�ӵ������������ݶ��롣"FALLING" - ���ʱ�ӵ��½��������ݶ���
	parameter	FVAL_LVAL_ALIGN			= "TRUE"				;	//"TRUE" - fval �� lval ֮��ľ���̶�Ϊ3��ʱ�ӡ�"FALSE" - fval �� lval ֮��ľ��������趨
	parameter	SOURCE_FILE_PATH		= "file/source_file/"	;	//����Դ�ļ�·��
	parameter	GEN_FILE_EN				= 0						;	//0-���ɵ�ͼ��д���ļ���1-���ɵ�ͼ��д���ļ�
	parameter	GEN_FILE_PATH			= "file/gen_file/"		;	//����������Ҫд���·��
	parameter	NOISE_EN				= 0						;	//0-������������1-��������

	//	-------------------------------------------------------------------------------------
	//	dut paramter
	//	-------------------------------------------------------------------------------------
	parameter	SENSOR_DAT_WIDTH		= 10	;	//sensor ���ݿ��
	parameter	REG_WD					= 32	;	//�Ĵ���λ��

	//	-------------------------------------------------------------------------------------
	//	monitor paramter
	//	-------------------------------------------------------------------------------------
	parameter	MONITOR_OUTPUT_FILE_EN			= 0						;	//�Ƿ��������ļ�
	parameter	MONITOR_OUTPUT_FILE_PATH		= "file/sync_buffer_file/"	;	//����������Ҫд���·��
	parameter	CHK_INOUT_DATA_STOP_ON_ERROR	= 0						;
	parameter	CHK_PULSE_WIDTH_STOP_ON_ERROR	= 0						;

	//	-------------------------------------------------------------------------------------
	//	testcase parameter
	//	-------------------------------------------------------------------------------------
	parameter	CLK_PERIOD				= 10	;	//ʱ��Ƶ�ʣ�100MHz

	//	===============================================================================================
	//	--ref signal
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	sensor signal
	//	-------------------------------------------------------------------------------------
	reg					clk_mt9p031		= 1'b0;
	reg					clk_pix			= 1'b0;
	wire				o_fval_mt9p031	;

	//	-------------------------------------------------------------------------------------
	//	dut signal
	//	-------------------------------------------------------------------------------------
	wire											o_fval_sensor	;
	wire											o_lval_sensor	;
	wire	[SENSOR_DAT_WIDTH*CHANNEL_NUM-1:0]		ov_pix_data_sensor	;
	wire											clk_sensor_pix	;
	wire											i_clk_en	;

	//	ref ARCHITECTURE

	//	===============================================================================================
	//	ref ***tb ��ģ�鼤��***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	--ref Sensor
	//	-------------------------------------------------------------------------------------
	always	#(CLK_PERIOD/2.0)	clk_mt9p031	= !clk_mt9p031;

	initial begin
		driver_mt9p031.bfm_mt9p031.reset_high();
		#200;
		driver_mt9p031.bfm_mt9p031.reset_low();
	end

	assign	o_fval_mt9p031	= harness.o_fval;

	//	-------------------------------------------------------------------------------------
	//	--ref DUT
	//	-------------------------------------------------------------------------------------
	always	#(CLK_PERIOD/2.0)		clk_pix		= !clk_pix;
	assign	o_fval_sensor			= driver_mt9p031.o_fval;
	assign	o_lval_sensor			= 1'b0;
	assign	ov_pix_data_sensor		= driver_mt9p031.ov_pix_data;
	assign	clk_sensor_pix			= driver_mt9p031.clk_sensor_pix;
	assign	i_clk_en				= 1'b1;

	//	-------------------------------------------------------------------------------------
	//	--ref ����ʱ��
	//	-------------------------------------------------------------------------------------
	initial begin
		#200
		//		repeat(20) @ (negedge harness.o_fval);
		repeat(30) @ (negedge driver_mt9p031.o_fval);
		#200
		$stop;
	end

	//	===============================================================================================
	//	ref ***����bfm task***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	--ref sensor pattern
	//	-------------------------------------------------------------------------------------
	//	initial begin
	//		forever begin
	//			driver_mt9p031.bfm_mt9p031.pattern_random(16,400);
	//		end
	//	end

	initial begin
		driver_mt9p031.bfm_mt9p031.pattern_2para(1,1);
	end

	//	-------------------------------------------------------------------------------------
	//	--ref ��ͣ��
	//	-------------------------------------------------------------------------------------
	initial begin
		harness.bfm_se_acq.acq_high();
		harness.bfm_se_acq.se_high();
		harness.bfm_reg_common.encrypt_high();
//		forever begin
//			harness.bfm_se_acq.se_acq_stop_start_random(1,2000);
//		end
	end

	initial begin
		forever begin
			harness.bfm_reg_common.pixel_format_random(20,1000);
		end
	end

	initial begin
		forever begin
			harness.bfm_reg_common.test_image_random(20,1000);
		end
	end
	
endmodule
