//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : harness
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/3/9 17:18:50	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------
`define		TESTCASE	testcase_1
module harness ();

	//	ref signals
	//	===============================================================================================
	//	--ref parameter
	//	===============================================================================================

	//	===============================================================================================
	//	--ref signal
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	����
	//	-------------------------------------------------------------------------------------
	wire								rst			;
	wire								wr_clk		;
	wire								rd_clk		;
	wire	[63:0]						din			;
	wire								wr_en		;
	wire								rd_en		;

	//	-------------------------------------------------------------------------------------
	//	���
	//	-------------------------------------------------------------------------------------
	wire	[31:0]						dout			;
	wire								full			;
	wire								empty			;
	wire								valid			;
	wire								prog_full		;
	wire								prog_empty		;


	//	ref ARCHITECTURE

	//	-------------------------------------------------------------------------------------
	//	���������ź�
	//	-------------------------------------------------------------------------------------
	assign	rst					= `TESTCASE.rst	;
	assign	wr_clk				= `TESTCASE.wr_clk	;
	assign	rd_clk				= `TESTCASE.rd_clk	;
	assign	din					= `TESTCASE.din	;
	assign	wr_en				= `TESTCASE.wr_en	;
	assign	rd_en				= `TESTCASE.rd_en	;



	//	-------------------------------------------------------------------------------------
	//	���� bfm ģ��
	//	-------------------------------------------------------------------------------------
	//	bfm_se_acq		bfm_se_acq();
	//
	//	bfm_reg_common # (
	//	.REG_WD		(`TESTCASE.REG_WD	)
	//	)
	//	bfm_reg_common ();


	//	-------------------------------------------------------------------------------------
	//	���� fifo ģ��
	//	-------------------------------------------------------------------------------------
	fifo_w64d256_pf180_pe6 fifo_w64d256_pf180_pe6_inst (
	.rst			(rst			),
	.wr_clk			(wr_clk			),
	.din			(din			),
	.wr_en			(wr_en			),
	.full			(full			),
	.prog_full		(prog_full		),
	.rd_clk			(rd_clk			),
	.rd_en			(rd_en			),
	.dout			(dout			),
	.empty			(empty			),
	.valid			(				),
	.prog_empty		(prog_empty		)
	);


	//generate vcd file
	//initial begin
	//$dumpfile("test.vcd");
	//$dumpvars(1,top_frame_buffer_inst);
	//end

	//for lattice simulation
	//GSR   GSR_INST (.GSR (1'b1)); //< global reset sig>
	//PUR   PUR_INST (.PUR (1'b1)); //<powerup reset sig>



endmodule
