//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : testcase_2
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/4/10 16:50:28	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ���ڴ�С��16x16�������ź���Ч������ģʽ�µ�����״��
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module testcase_2 ();

	//	ref signals
	//	===============================================================================================
	//	--ref parameter
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	TESTCASE
	//	-------------------------------------------------------------------------------------
	parameter	TESTCASE_NUM			= "testcase_2"			;	//����ģ����Ҫʹ���ַ���
	//	-------------------------------------------------------------------------------------
	//	dut paramter
	//	-------------------------------------------------------------------------------------
	parameter	FIFO_WIDTH		= 8		;
	parameter	FIFO_DEPTH		= 16	;

	//	-------------------------------------------------------------------------------------
	//	monitor paramter
	//	-------------------------------------------------------------------------------------
	parameter	MONITOR_OUTPUT_FILE_EN			= 0						;	//�Ƿ��������ļ�
	parameter	MONITOR_OUTPUT_FILE_PATH		= "file/sync_buffer_file/"	;	//����������Ҫд���·��
	parameter	CHK_INOUT_DATA_STOP_ON_ERROR	= 0						;
	parameter	CHK_PULSE_WIDTH_STOP_ON_ERROR	= 0						;

	//	-------------------------------------------------------------------------------------
	//	testcase parameter
	//	-------------------------------------------------------------------------------------
	parameter	CLK_PERIOD_WR				= 15	;	//ʱ��Ƶ��
	parameter	CLK_PERIOD_RD				= 23	;	//ʱ��Ƶ��

	//	===============================================================================================
	//	--ref signal
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	dut signal
	//	-------------------------------------------------------------------------------------
	reg								reset_async		= 1'b0	;
	reg								clk_wr			= 1'b0	;
	reg								i_wr_en			= 1'b0	;
	reg		[FIFO_WIDTH-1:0]		iv_fifo_din		= 'b0	;
	reg								clk_rd			= 1'b0	;
//	wire							i_rd_en			;
	reg								i_rd_en			= 1'b0	;

	//	-------------------------------------------------------------------------------------
	//	testbench
	//	-------------------------------------------------------------------------------------
	reg								rd_begin		= 1'b0;

	//	ref ARCHITECTURE

	//	===============================================================================================
	//	ref ***tb ��ģ�鼤��***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	--ref DUT
	//	-------------------------------------------------------------------------------------
	//	-------------------------------------------------------------------------------------
	//	ʱ�Ӹ�λ
	//	-------------------------------------------------------------------------------------
	always	#(CLK_PERIOD_WR/2.0)	clk_wr	= !clk_wr;
	always	#(CLK_PERIOD_RD/2.0)	clk_rd	= !clk_rd;

	initial begin
		reset_async	= 1'b1;
		#200;
		reset_async	= 1'b0;
	end

	//	-------------------------------------------------------------------------------------
	//	д
	//	-------------------------------------------------------------------------------------
	//	always @ (posedge clk_wr) begin
	//		i_wr_en	<= $random();
	//	end

	initial begin
		forever begin
			wait(harness.o_fifo_full==1'b0 && harness.o_fifo_empty==1'b1);
			@(posedge clk_wr);
			i_wr_en	= 1'b1;
			wait(harness.o_fifo_full==1'b1);
			@(posedge clk_wr);
			i_wr_en	= 1'b0;
		end
	end

	always @ (posedge clk_wr) begin
		if((i_wr_en==1)&&(harness.o_fifo_full==1'b0)) begin
			iv_fifo_din	<= iv_fifo_din + 1'b1;
		end
	end

	//	-------------------------------------------------------------------------------------
	//	��
	//	-------------------------------------------------------------------------------------
	initial begin
		forever begin
			wait(harness.o_fifo_full==1'b1 && harness.o_fifo_empty==1'b0);
			@(posedge clk_rd);
			i_rd_en	= 1'b1;
			wait(harness.o_fifo_empty==1'b1);
			@(posedge clk_rd);
			i_rd_en	= 1'b0;
		end
	end

	//	-------------------------------------------------------------------------------------
	//	--ref ����ʱ��
	//	-------------------------------------------------------------------------------------
	initial begin
		#200
		#10000
		#200
		$stop;
	end


endmodule
