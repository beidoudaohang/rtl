
//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : ccd_count.v
//  -- �����       : ��
//-------------------------------------------------------------------------------------------------
//
//  --�޸ļ�¼  :
//
//  -- ����         :| �޸�����     :|  �޸�˵��
//---------------------------------------------------------------------------------------
//  -- ��       	:| 09/01/2013   :|  ��ʼ�汾
//  -- ��Сƽ      	:| 04/29/2015   :|  �����޸ģ���Ӧ��ICX445 sensor
//  -- �Ϻ���      	:| 2015/12/8    :|  ��ֲ��u3
//---------------------------------------------------------------------------------------
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ����CCD������
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale      1ns/100ps
//-------------------------------------------------------------------------------------------------

module ccd_count # (
	parameter	LINE_PERIOD		= 1532		,	//������
	parameter	LINE_CNT_WIDTH	= 13			//�м��������
	)
	(
	input							clk     	,   //ʱ��
	input							reset		,	//
	output							o_line_end	,	//
	output	[LINE_CNT_WIDTH-1:0]	ov_count		//
	);

	//	ref signals
	//	-------------------------------------------------------------------------------------
	//	�źŶ���
	//	-------------------------------------------------------------------------------------
	reg		[LINE_CNT_WIDTH-1:0]		count		= 'b0;
	reg									line_end	= 1'b0;

	//	ref ARCHITECTURE
	//  ===============================================================================================
	//  �ڶ����֣��������߼�
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//  ����˵�����������ڼ�����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(reset) begin
			count	<= 'b0;
		end
		else if(count==(LINE_PERIOD-1)) begin
			count	<= 'b0;
		end
		else begin
			count	<= count + 1'b1;
		end
	end
	assign	ov_count	= count;

	//  -------------------------------------------------------------------------------------
	//  ����˵�����������ڱ�־
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(count==(LINE_PERIOD-2)) begin
			line_end	<= 1'b1;
		end
		else begin
			line_end	<= 1'b0;
		end
	end
	assign	o_line_end	= line_end;

endmodule