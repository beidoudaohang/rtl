//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : fifo_con
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2013/6/13 10:17:01	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :	ǰ��FIFO�ĸ�λģ�飬����1CLK�ĸ�λ�ź�
//              1)  : �첽FIFO�Ķ�д�˿���Ҫ�Ը�λ�ź�ͬ����������ڸ���ʱ�����3�������ڣ�FIFO���ǳ��ڸ�λ״̬
//
//              2)  : fval��dval֮��Ҫ���㹻�Ŀ�϶
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//`include			"frame_buffer_def.v"
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module fifo_con (
	input			clk			,
	input			i_fval		,
	output			o_rst_buf
	);

	//ref signals
	reg				fval_d 		= 1'b0;
	reg				buf_rst_reg = 1'b0;
	wire			fval_rise	;

	//ref ARCHITECTURE

	//��fval�����ص���ʱ����λǰ��FIFO
	always @ (posedge clk) begin
		fval_d		<= i_fval;
		buf_rst_reg	<= fval_rise;
	end

	assign	fval_rise	= (~fval_d)&i_fval;
	assign	o_rst_buf	= buf_rst_reg;


endmodule
