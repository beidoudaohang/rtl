//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : wb_statis
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/2/13 10:30:32	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ����ǰ�������ͳ��������ɷ���ͳ��
//              1)  : G����ͳ��ֵ/2 ��������ͳ��ֵ����
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module wb_statis # (
	parameter					SENSOR_DAT_WIDTH	= 10	,	//sensor ���ݿ��
	parameter					WB_STATIS_WIDTH		= 29	,	//��ƽ��ģ��ͳ��ֵ���
	parameter					REG_WD				= 32		//�Ĵ���λ��
	)
	(
	input							clk						,	//����ʱ��
	input							i_fval					,	//���ź�
	input							i_lval					,	//���ź�
	input	[SENSOR_DAT_WIDTH-1:0]	iv_pix_data				,	//ͼ������
	input							i_r_flag				,	//��ɫ������־ R
	input							i_g_flag				,	//��ɫ������־ G
	input							i_b_flag				,	//��ɫ������־ B
	input							i_interrupt_pin			,	//�ж�ģ��������ж��źţ�1-�ж���Ч�����ж�������ʱ��������ɫ����ͳ��ֵ�ʹ��ڼĴ������˿�
	output	[WB_STATIS_WIDTH-1:0]	ov_wb_statis_r			,	//������ظ�ʽΪ8bit����ֵΪͼ��R����8bitͳ��ֵ��������ظ�ʽΪ����8bit����ֵΪͼ��R������8bitͳ��ֵ��
	output	[WB_STATIS_WIDTH-1:0]	ov_wb_statis_g			,	//������ظ�ʽΪ8bit����ֵΪͼ��G����8bitͳ��ֵ����2�Ľ����������ظ�ʽΪ����8bit����ֵΪͼ��G������8bitͳ��ֵ����2�Ľ����
	output	[WB_STATIS_WIDTH-1:0]	ov_wb_statis_b				//������ظ�ʽΪ8bit����ֵΪͼ��B����8bitͳ��ֵ��������ظ�ʽΪ����8bit����ֵΪͼ��B������8bitͳ��ֵ��
	);

	//	ref signals

	reg								fval_dly0			= 1'b0;
	reg								fval_dly1			= 1'b0;
	wire							fval_rise			;
	reg								int_pin_dly			= 1'b0;
	wire							int_pin_rise		;
	reg		[WB_STATIS_WIDTH-1:0]	wb_statis_r			= {WB_STATIS_WIDTH{1'b0}};
	reg		[WB_STATIS_WIDTH:0]		wb_statis_g			= {(WB_STATIS_WIDTH+1){1'b0}};
	reg		[WB_STATIS_WIDTH-1:0]	wb_statis_b			= {WB_STATIS_WIDTH{1'b0}};
	reg		[WB_STATIS_WIDTH-1:0]	wb_statis_r_reg		= {WB_STATIS_WIDTH{1'b0}};
	reg		[WB_STATIS_WIDTH-1:0]	wb_statis_g_reg		= {WB_STATIS_WIDTH{1'b0}};
	reg		[WB_STATIS_WIDTH-1:0]	wb_statis_b_reg		= {WB_STATIS_WIDTH{1'b0}};


	//	ref ARCHITECTURE

	//  ===============================================================================================
	//	ref ***��ʱ ȡ����***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	����Чȡ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_dly0	<= i_fval;
	end
	assign	fval_rise	= (fval_dly0==1'b0 && i_fval==1'b1) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//	�ж�ȡ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		int_pin_dly	<= i_interrupt_pin;
	end
	assign	int_pin_rise	= (int_pin_dly==1'b0 && i_interrupt_pin==1'b1) ? 1'b1 : 1'b0;

	//  ===============================================================================================
	//	ref ***ͳ����ɫ����***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	r����
	//	1.����������ʱ����λ�ڲ�������
	//	2.��������־��Чʱ�������������������
	//	3.��ɫ������־ֻ��lval��Чʱ=1����˲���Ҫlval��Ϊ����
	//	4.ֻͳ�Ƹ�8bit
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(fval_rise) begin
			wb_statis_r	<= {WB_STATIS_WIDTH{1'b0}};
		end
		else begin
			if(i_r_flag) begin
				wb_statis_r	<= wb_statis_r + iv_pix_data[SENSOR_DAT_WIDTH-1:SENSOR_DAT_WIDTH-8];
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	g����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(fval_rise) begin
			wb_statis_g	<= {(WB_STATIS_WIDTH+1){1'b0}};
		end
		else begin
			if(i_g_flag) begin
				wb_statis_g	<= wb_statis_g + iv_pix_data[SENSOR_DAT_WIDTH-1:SENSOR_DAT_WIDTH-8];
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	g����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(fval_rise) begin
			wb_statis_b	<= {WB_STATIS_WIDTH{1'b0}};
		end
		else begin
			if(i_b_flag) begin
				wb_statis_b	<= wb_statis_b + iv_pix_data[SENSOR_DAT_WIDTH-1:SENSOR_DAT_WIDTH-8];
			end
		end
	end

	//  ===============================================================================================
	//	ref ***���ͳ�ƽ��***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	r���������ж��źŵ������أ����ڲ�ͳ�ƽ�����浽�˿���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(int_pin_rise) begin
			wb_statis_r_reg	<= wb_statis_r;
		end
	end
	assign	ov_wb_statis_r	= wb_statis_r_reg;

	//  -------------------------------------------------------------------------------------
	//	g���������ж��źŵ������أ����ڲ�ͳ�ƽ�����浽�˿��ϣ����ֵҪ����2
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(int_pin_rise) begin
			wb_statis_g_reg	<= wb_statis_g[WB_STATIS_WIDTH:1];
		end
	end
	assign	ov_wb_statis_g	= wb_statis_g_reg;

	//  -------------------------------------------------------------------------------------
	//	b���������ж��źŵ������أ����ڲ�ͳ�ƽ�����浽�˿���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(int_pin_rise) begin
			wb_statis_b_reg	<= wb_statis_b;
		end
	end
	assign	ov_wb_statis_b	= wb_statis_b_reg;


endmodule