//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : leader
//  -- �����       : ��ǿ
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- ��ǿ         :| 2014/12/3 13:58:33	:|  ���ݼ���Ԥ������
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������
//              1)  : U3V��ʽleaderģ�飬��ϳɷ���U3V��ʽleader��
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------
module leader #(
	parameter							DATA_WD			= 32	,	//�����������λ������ʹ��ͬһ���
	parameter							SHORT_REG_WD	= 16	,	//�̼Ĵ���λ��
	parameter							REG_WD 			= 32	,	//�Ĵ���λ��
	parameter							LONG_REG_WD 	= 64		//���Ĵ���λ��
	)
	(
//  ===============================================================================================
//  ��һ���֣�ʱ�Ӹ�λ
//  ===============================================================================================
	input								reset					,		//��λ�źţ��ߵ�ƽ��Ч������ʱ��ʱ����
	input								clk						,		//ʱ���źţ�����ʱ��ʱ����ͬ�ڲ�����ʱ��
//  ===============================================================================================
//  �ڶ����֣�ͷ����־
//  ===============================================================================================
	input								i_leader_flag			,		//ͷ����־
//  ===============================================================================================
//  �������֣����ƼĴ�����chunk��Ϣ��ֻ���Ĵ���
//  ===============================================================================================
	input		[REG_WD-1			:0]	iv_pixel_format         ,       //���ظ�ʽ�����������leader��
	input								i_chunk_mode_active     ,       //chunk�ܿ��أ����ش�Payload Typeʹ��Ϊimage extend chunk ���ͣ�chunk�ر�Ϊimage����
	input		[LONG_REG_WD-1		:0]	iv_blockid				,		//ͷ����chunk��β����blockid��Ϣ����һ֡��block ID��0��ʼ��������һ֡block IDΪ0
	input		[LONG_REG_WD-1		:0]	iv_timestamp			, 		//ͷ���е�ʱ����ֶ�,iv_timestamp�ڳ��ź�������8��ʱ��֮������ȶ�
	input		[SHORT_REG_WD-1		:0]	iv_size_x				, 		//ͷ���еĴ��ڿ��
	input		[SHORT_REG_WD-1		:0]	iv_size_y				, 		//ͷ���еĴ��ڸ߶�
	input		[SHORT_REG_WD-1		:0]	iv_offset_x				, 		//ͷ���е�ˮƽƫ��
	input		[SHORT_REG_WD-1		:0]	iv_offset_y				, 		//ͷ���еĴ�ֱ����

//  ===============================================================================================
//  ���Ĳ��֣�������Ч������
//  ===============================================================================================
	output	reg							o_data_valid			,       //�����ͷ��������Ч�ź�
	output	reg	[DATA_WD-1			:0]	ov_data                         //ͷ������
	);
//  ===============================================================================================
//  ���ز���
//  ===============================================================================================
	localparam							LEADER_LENTH	=	4'd13	;		//ͷ������13
//  ===============================================================================================
//  �����ͼĴ�������
//  ===============================================================================================
	reg			[3					:0]	count          = 	4'h0;		//���������������ͷ���е��ź�
//  ===============================================================================================
//  i_leader_flag�ڼ���
//  ===============================================================================================
	always @ (posedge clk) begin
		if(i_leader_flag) begin
			count	<=	count + 4'h1;
		end
		else begin
			count	<=	4'h0;
		end
	end
//  -------------------------------------------------------------------------------------
//  ����leader�����ݣ�����ʽ����Image Extended Chunk Leader��ʽ
//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if ( reset ) begin
			ov_data <= 	32'h0;
		end
		else  begin
			case ( count )
				4'h1	:	ov_data	<=	32'h4c563355				;
				4'h2	:   ov_data	<=	{16'd52,16'd0}				;
				4'h3	:   ov_data	<=	iv_blockid[31:0]          	;
				4'h4	:   ov_data	<=	iv_blockid[63:32]         	;
				4'h5	:   ov_data	<=	{1'b0,i_chunk_mode_active,{14'h0001},16'h0000}	;	//����ֻ֧��Image��0x0001����Image Extended Chunk��0x4001��
				4'h6	:   ov_data	<=	iv_timestamp[31:0]			;
				4'h7	:   ov_data	<=	iv_timestamp[63:32]			;
				4'h8	:   ov_data	<=	iv_pixel_format				;
				4'h9	:   ov_data	<=	{16'h00,iv_size_x}			;
				4'ha	:   ov_data	<=	{16'h00,iv_size_y}			;
				4'hb	:   ov_data	<=	{16'h00,iv_offset_x}		;
				4'hc	:   ov_data	<=	{16'h00,iv_offset_y}		;
				4'hd	:   ov_data	<=	32'h0						;
				default	:  	ov_data <= 	32'h0						;
			endcase
		end
	end
//  -------------------------------------------------------------------------------------
//  ���o_data_valid�ź�
//  -------------------------------------------------------------------------------------
	always @ (posedge clk ) begin
		if ( reset ) begin
			o_data_valid	<=	1'b0;
		end
		else if (( count>4'h0 ) && ( count <= LEADER_LENTH ))begin
			o_data_valid	<=	1'b1;
		end
		else begin
			o_data_valid	<=	1'b0;
		end
	end

endmodule