//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : ad_output_latch
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/8/9 14:16:15	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module ad_output_latch (
	input				clk					,	//����ʱ��
	input	[13:0]		iv_pix_data			,	//��������
	input				i_lvds_pattern_en	,	//lvds������ʹ��
	input	[15:0]		iv_lvds_pattern		,	//lvds������
	input				i_sync_word_sel		,	//ͬ����ѡ���ź�
	input	[15:0]		iv_sync_word		,	//ͬ����
	output	[15:0]		ov_pix_data				//�����������
	);

	//	ref signals
	reg		[15:0]			pattern_mux		= 16'b0;
	reg		[15:0]			pattern_mux_dly	= 16'b0;
	reg		[15:0]			pix_data_reg	= 16'b0;


	//	ref ARCHITECTURE

	//	-------------------------------------------------------------------------------------
	//	������ѡ��mux
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(i_lvds_pattern_en) begin
			pattern_mux	<= iv_lvds_pattern;
		end
		else begin
			pattern_mux	<= {iv_pix_data,2'b00};
		end
	end

	//	-------------------------------------------------------------------------------------
	//	��ʱ1��
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		pattern_mux_dly	<= pattern_mux;
	end

	//	-------------------------------------------------------------------------------------
	//	�滻ͬ����
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(i_sync_word_sel) begin
			pix_data_reg	<= iv_sync_word;
		end
		else begin
			pix_data_reg	<= pattern_mux_dly;
		end
	end
	assign	ov_pix_data	= pix_data_reg	;



endmodule
