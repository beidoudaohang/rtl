
//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : ccd_exp.v
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  --�޸ļ�¼  :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���      	:| 2015/12/23 10:51:52	:|  ��ʼ�汾����mv_ccd���޸�
//-------------------------------------------------------------------------------------------------
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ccd_exp �����ع���ֱ�־
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale      1ns/100ps
//-------------------------------------------------------------------------------------------------

module ccd_exp # (
	parameter	LINE_PERIOD		= 1532		,	//������
	parameter	LINE_CNT_WIDTH	= 13			//�м��������
	)
	(
	input									clk      			,   //ʱ��
	input									reset				,	//��λ������Ч
	input		[`EXP_WD-1:0]				iv_exp_reg			,   //�ع�ʱ�Ӹ����Ĵ���
	input		[`EXP_WD-1:0]				iv_exp_line_reg		,	//�ع�����ʱ�Ӹ����Ĵ���
	input		[`FRAME_WD-1:0]				iv_exp_start_reg	,	//
	input  		[`FRAME_WD-1:0]				iv_vcount			,	//
	input									i_readout_flag		,	//
	input                       			i_start_acquisit	,   //��CCDģ��Ŀ����ź�
	input									i_triggermode		,   //��CCDģ��Ĳɼ�ģʽ�ź�
	input									i_trigger			,   //��CCDģ��Ĵ����ź�
	input									i_xsg_flag			,	//
	input									i_exposure_end		,	//
	output									o_reg_active		,	//
	output		[LINE_CNT_WIDTH-1:0]		ov_hcount			,	//�м�����
	output  								o_line_end			,	//�н�����־�����м����������ֵ����
	output									o_exp_line_end		,	//�ع��н�����־
	output									o_trigger_mask		,	//���α�־
	output									o_integration       	//�����ź�
	);

	//	ref signals
	wire							hcount_reset				;
	reg			[3:0]				start_acquisit_shift		;
	reg			[1:0]				triggermode_shift			;
	reg			[1:0]				exp_start_line_flag_shift	;
	wire							exp_start_line_flag			;
	reg								trigger_reg					;
	reg								trigger_reg_dly_0			;
	reg								trigger_reg_dly_1			;
	reg								trigger2hend				;
	wire							exp_start_tri				;
	wire							exp_start_con				;
	wire							exp_start					;
	reg								exp_flag 					;
	reg		[`EXP_WD-1:0]			exp_count					;
	wire							integration_start			;
	reg								trig_2_cont_wt_hend			;
	reg		[1:0]					xsg_flag_shift				;

	//	ref ARCHITECTURE

	//  ===============================================================================================
	//  �ڶ����֣�ģ��ʵ����
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//  ccd_count		: ccd���ڼ�����
	//  -------------------------------------------------------------------------------------
	ccd_count # (
	.LINE_PERIOD	(LINE_PERIOD	),
	.LINE_CNT_WIDTH	(LINE_CNT_WIDTH	)
	)
	ccd_count_inst (
	.clk			(clk			),
	.reset			(hcount_reset	),
	.o_line_end		(o_line_end		),
	.ov_count		(ov_hcount		)
	);

	//  ===============================================================================================
	//  �������֣��ع���ʼ�߼�
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	i_start_acquisit ȡ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		start_acquisit_shift	<= {start_acquisit_shift[2:0],i_start_acquisit};
	end

	//  -------------------------------------------------------------------------------------
	//	i_triggermode ȡ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		triggermode_shift	<= {triggermode_shift[0],i_triggermode};
	end

	//  -------------------------------------------------------------------------------------
	//	exp_start_line_flag ȡ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		exp_start_line_flag_shift	<= {exp_start_line_flag_shift[0],exp_start_line_flag};
	end

	//  -------------------------------------------------------------------------------------
	//	����˵���������ع⿪ʼ�б�־
	//  -------------------------------------------------------------------------------------
	assign exp_start_line_flag	= (iv_exp_start_reg==iv_vcount) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//  ����ģʽ�ع�����ν׶�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(reset) begin
			trigger_reg	<= 1'b0;
		end
		else if(!o_trigger_mask && i_triggermode && i_start_acquisit) begin
			trigger_reg <= i_trigger;
		end
		else begin
			trigger_reg	<= 1'b0;
		end
	end

	always @ (posedge clk) begin
		trigger_reg_dly_0	<= trigger_reg;
		trigger_reg_dly_1	<= trigger_reg_dly_0;
	end

	//  -------------------------------------------------------------------------------------
	//  ����ģʽ�عⷢ����i_readout_flag��Чʱ,������hend
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(reset) begin
			trigger2hend	<=	1'b0;
		end
		else if(trigger_reg_dly_1 && i_readout_flag) begin
			trigger2hend	<=	1'b1;
		end
		else if(o_line_end) begin
			trigger2hend	<=	1'b0;
		end
	end

	//  -------------------------------------------------------------------------------------
	// ����������ʱ����readout�׶Σ�,������hend������һ�п�ʼ�������ع�
	//  -------------------------------------------------------------------------------------

	always @ ( posedge clk )
	begin
		if(reset)
		begin
			trig_2_cont_wt_hend	<=	1'b0;
		end
		else if((triggermode_shift == 2'b10) && !o_trigger_mask)
		begin
			trig_2_cont_wt_hend	<=	1'b1;
		end
		else if(o_line_end)
		begin
			trig_2_cont_wt_hend	<=	1'b0;
		end
	end
	//  -------------------------------------------------------------------------------------
	//  ���ֲ�ͬ�ع�ģʽ��ʼ�ź�
	//	����ģʽʱ��1������������
	//				2�������ع���ʼ�б�־
	//
	//	����ģʽʱ��1�������Ҵ������ع�����ν׶�
	//
	//	����ģʽ�л�������ģʽ��!i_readout_flagʱ
	//		����������ʱ�������ν׶Σ������ع���ʼ�׶Σ��ӳٵ���hendʱ���ٿ�ʼ�ع⣨��Сƽ����
	//  -------------------------------------------------------------------------------------

	assign	exp_start_tri 	= (trigger2hend && o_line_end) || (trigger_reg_dly_1 && !i_readout_flag)											;
	assign	exp_start_con 	= ((start_acquisit_shift == 4'b0111) || (exp_start_line_flag && o_line_end)) || (trig_2_cont_wt_hend & o_line_end)		;
	assign	exp_start 		= i_start_acquisit ? (i_triggermode ? exp_start_tri : exp_start_con) : 1'b0										;

	//  -------------------------------------------------------------------------------------
	//  ����˵����w_hcount_set
	//	����������
	//		1���عⷢ����i_readout_flag��Чʱ	��	��λhcount
	//  -------------------------------------------------------------------------------------
	assign	hcount_reset 	= (!i_readout_flag & exp_start) ;

	//  ===============================================================================================
	//  ���Ĳ��֣������ع������
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//  ����˵���������ع����ڼ�������������ʱ��Ϊ��λ
	//  -------------------------------------------------------------------------------------

	always @ ( posedge clk )
	begin
		if(reset)
		begin
			exp_flag	<=	1'b0;
		end
		else if((exp_count == iv_exp_reg) || !i_start_acquisit)
		begin
			exp_flag	<=	1'b0;
		end
		else if(exp_start)
		begin
			exp_flag	<=	1'b1;
		end
	end

	always @ ( posedge clk )
	begin
		if(reset)
		begin
			exp_count	<=	`EXP_WD'h0;
		end
		else if(exp_flag)
		begin
			exp_count	<=	exp_count + `EXP_WD'h1;
		end
		else
		begin
			exp_count	<=	`EXP_WD'h0;
		end
	end

	//  ===============================================================================================
	//  ���岿�֣�����ع���ر�־
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//  ����˵���� �ع�����
	//  -------------------------------------------------------------------------------------

	assign	integration_start	= ((exp_count == `SUB_PER_WIDTH) && exp_flag && i_start_acquisit) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//  ����˵���� ���ع����������XSG�׶�
	//  -------------------------------------------------------------------------------------

	assign	o_exp_line_end		= ((exp_count == iv_exp_line_reg) && exp_flag && i_start_acquisit) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//  ����˵�������ֱ�־
	//  -------------------------------------------------------------------------------------

	always @ ( posedge clk )
	begin
		if(reset)
		begin
			o_integration	<= 1'b0;
		end
		else if(i_exposure_end || !i_start_acquisit)
		begin
			o_integration 	<= 1'b0;
		end
		else if(integration_start)
		begin
			o_integration 	<= 1'b1;
		end
	end

	//  -------------------------------------------------------------------------------------
	//  ����˵�����ع����α�־
	//  -------------------------------------------------------------------------------------

	always @ ( posedge clk )
	begin
		if(reset)
		begin
			o_trigger_mask	<= 1'b0;
		end
		else if((exp_start_line_flag_shift == 2'b01) || !i_start_acquisit)
		begin
			o_trigger_mask 	<= 1'b0;
		end
		else if(exp_start || trigger_reg)
		begin
			o_trigger_mask 	<= 1'b1;
		end
	end

	//  ===============================================================================================
	//  �������֣��Ĵ�����Чʱ��
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	xsg_flag_shift ȡ��
	//  -------------------------------------------------------------------------------------

	always @ ( posedge clk )
	begin
		xsg_flag_shift	<=	{xsg_flag_shift[0],i_xsg_flag};
	end

	//  -------------------------------------------------------------------------------------
	//	����˵����
	//		1������ģʽ�¿���ʱ
	//		2���ع������ʼ�µĴ���֡ʱ
	//		3������ģʽʱ����������֡���ٴ���ʱ
	//  -------------------------------------------------------------------------------------

	assign	o_reg_active =  (start_acquisit_shift == 4'b0001) || (i_triggermode && !i_readout_flag && trigger_reg) || (xsg_flag_shift == 2'b10);

endmodule