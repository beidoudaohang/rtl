//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : grey_statis
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/3/18 15:16:24	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : �Ҷ�ͳ��ģ��
//              1)  : ���� aoi �г��źţ��ۼ�ÿ������
//
//              2)  : o_fval��ʱ1��ʱ��
//
//              3)  : ���ظ�ʽ8bit-ͳ�Ƶ�8bit������-ȫ��ͳ��
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module grey_statis # (
	parameter						SENSOR_DAT_WIDTH	= 10	,	//sensor ���ݿ��
	parameter						GREY_STATIS_WIDTH	= 48	,	//�Ҷ�ͳ��ģ��ͳ��ֵ���
	parameter						REG_WD				= 32		//�Ĵ���λ��
	)
	(
	//Sensor�����ź�
	input								clk						,	//����ʱ��
	input								i_fval					,	//���ź�
	input								i_lval					,	//���ź�
	input	[SENSOR_DAT_WIDTH-1:0]		iv_pix_data				,	//ͼ������
	//����ģ������
	input								i_interrupt_pin			,	//�ж�ģ��������ж��źţ�1-�ж���Ч�����ж�������ʱ������Ҷ�ͳ��ֵ�ʹ��ڼĴ������˿�
	//�Ҷ�ͳ����ؼĴ���
	input	[REG_WD-1:0]				iv_pixel_format			,	//���ظ�ʽ�Ĵ���0x01080001:Mono8��0x01100003:Mono10��0x01080008:BayerGR8��0x0110000C:BayerGR10
	output	[GREY_STATIS_WIDTH-1:0]		ov_grey_statis_sum			//�üĴ���ֵΪͼ��Ҷ�ͳ��ֵ�ܺ͡�������ظ�ʽΪ8bit����ֵΪ����8bitͳ��ֵ��������ظ�ʽΪ10bit����ֵΪ����10bitͳ��ֵ
	);

	//	ref signals

	reg									fval_dly0		= 1'b0;
	reg									fval_dly1		= 1'b0;
	wire								fval_rise		;
	reg									int_pin_dly		= 1'b0;
	wire								int_pin_rise	;
//	reg									format8_sel		= 1'b0;
	reg		[GREY_STATIS_WIDTH-1:0]		grey_statis		= {GREY_STATIS_WIDTH{1'b0}};
	reg		[GREY_STATIS_WIDTH-1:0]		grey_statis_reg	= {GREY_STATIS_WIDTH{1'b0}};



	//	ref ARCHITECTURE


	//  ===============================================================================================
	//	ref ***��ʱ ȡ����***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	����Чȡ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_dly0	<= i_fval;
	end
	assign	fval_rise	= (fval_dly0==1'b0 && i_fval==1'b1) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//	�ж�ȡ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		int_pin_dly	<= i_interrupt_pin;
	end
	assign	int_pin_rise	= (int_pin_dly==1'b0 && i_interrupt_pin==1'b1) ? 1'b1 : 1'b0;

	//  ===============================================================================================
	//	ref ***ͳ������***
	//  ===============================================================================================
	//	//  -------------------------------------------------------------------------------------
	//	//	Mono8		- 0x01080001	-> 0x1081	-> 0001,0000,1000,,,,0001
	//	//	Mono10		- 0x01100003	-> 0x1103	-> 0001,0001,0000,,,,0011
	//	//	BayerGR8	- 0x01080008	-> 0x1088	-> 0001,0000,1000,,,,1000
	//	//	BayerGR10	- 0x0110000C	-> 0x110C	-> 0001,0001,0000,,,,1100
	//	//											   --------!-!-------!!!!
	//	//                                                     ^    ^       ^------bit0
	//	//                                             bit20---|    |---bit16
	//	//	����� ! �ģ����ǲ���Ƚϵ�bit.�ֱ��� bit
	//	//  -------------------------------------------------------------------------------------
	//	//  -------------------------------------------------------------------------------------
	//	//	format8_sel
	//	//	1.�ж����ظ�ʽ�Ƿ�ѡ��8bit���ظ�ʽ
	//	//	2.ʹ��6bit�ж�����
	//	//  -------------------------------------------------------------------------------------
	//	always @ (posedge clk) begin
	//		case({iv_pixel_format[20],iv_pixel_format[19],iv_pixel_format[3:0]})
	//			6'b010001	: format8_sel	<= 1'b1;
	//			6'b011000	: format8_sel	<= 1'b1;
	//			default		: format8_sel	<= 1'b0;
	//		endcase
	//	end

	//	//  -------------------------------------------------------------------------------------
	//	//	�Ҷ�ͳ��ֵ
	//	//	1.����������ʱ����λ�ڲ�������
	//	//	2.lval��Чʱ�������������������
	//	//	3.���ظ�ʽ��8bitʱ��ͳ�Ƹ�8bit�����ظ�ʽ��10bit��ͳ��10bit��
	//	//  -------------------------------------------------------------------------------------
	//	always @ (posedge clk) begin
	//		if(fval_rise) begin
	//			grey_statis	<= {GREY_STATIS_WIDTH{1'b0}};
	//		end
	//		else begin
	//			if(i_lval) begin
	//				if(format8_sel) begin
	//					grey_statis	<= grey_statis + iv_pix_data[SENSOR_DAT_WIDTH-1:SENSOR_DAT_WIDTH-8];
	//				end
	//				else begin
	//					grey_statis	<= grey_statis + iv_pix_data[SENSOR_DAT_WIDTH-1:0];
	//				end
	//
	//			end
	//		end
	//	end

	//  -------------------------------------------------------------------------------------
	//	�Ҷ�ͳ��ֵ
	//	1.����������ʱ����λ�ڲ�������
	//	2.lval��Чʱ�������������������
	//	3.���ظ�ʽ��8bitʱ��ͳ��8bit�����ظ�ʽ��10bit��ͳ�Ƹ�8bit��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(fval_rise) begin
			grey_statis	<= {GREY_STATIS_WIDTH{1'b0}};
		end
		else begin
			if(i_lval) begin
				grey_statis	<= grey_statis + iv_pix_data[SENSOR_DAT_WIDTH-1:SENSOR_DAT_WIDTH-8];
			end
		end
	end

	//  ===============================================================================================
	//	ref ***���ͳ�ƽ��***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	���ж��źŵ������أ����ڲ�ͳ�ƽ�����浽�˿���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(int_pin_rise) begin
			grey_statis_reg	<= grey_statis;
		end
	end
	assign	ov_grey_statis_sum	= grey_statis_reg;


endmodule
