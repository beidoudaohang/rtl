//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : data_mask
//  -- �����       : �ܽ�
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �ܽ�       :| 2015/10/26 14:09:17	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : �������ɼ�ģʽ�£�ͨ�����е�ͼ������ݣ��ڴ����ɼ�ģʽ�£�ֻͨ��
//					����֡�����˳�����֮֡���ͼ�����ݡ�
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module data_mask #(
	parameter		SENSOR_DAT_WIDTH			= 12					,	//sensor ���ݿ��
	parameter		CHANNEL_NUM					= 4						,	//��������ͨ������
	parameter		CLK_FREQ_KHZ				= 55000					,	//ʱ��Ƶ�ʣ�55000KHz
	parameter		TRIGGER_STATUS_INTERVAL		= 1100					 	//trigger_status�쳣ʱ�䣬110ms
	)
	(
	input											clk					,	//ʱ��
	//�����ź�
	input											i_pll_lock			,	//�⴮ʱ���򣬽⴮pll�����ź�
	input											i_acquisition_start	,	//�����źţ�0-ͣ�ɣ�1-����
	input											i_stream_enable		,	//��ʹ���ź�
	input											i_trigger_start		,	//clk_pixʱ���򣬳������13��i2c��������.1:i2c restart���ʼ
	input											i_trigger_mode		,	//clk_pixʱ����ctrl_channel�����0-�����ɼ���1-�����ɼ�
	//ͼ������
	input											i_fval				,	//�⴮ʱ�������볡�ź�
	input											i_lval				,	//�⴮ʱ�����������ź�
	input	[SENSOR_DAT_WIDTH*CHANNEL_NUM-1:0]		iv_pix_data			,	//�⴮ʱ��������ͼ������
	//���trigger_mode�ź�
	output											o_trigger_mode		,	//�⴮ʱ�������trigger_mode�ź�
	output											o_trigger_status	,	//�⴮ʱ����1-�д����ź��Ҵ���֡δ�����ϣ�0-�޴����źŻ򴥷�֡������
	//����ź�
	output											o_fval				,	//�⴮ʱ����������ź�
	output											o_lval				,	//�⴮ʱ����������ź�
	output	[SENSOR_DAT_WIDTH*CHANNEL_NUM-1:0]		ov_pix_data			 	//�⴮ʱ�������ͼ������
	);

	//	ref signals


	//  -------------------------------------------------------------------------------------
	//	ref localparam
	//  -------------------------------------------------------------------------------------
	localparam	TRIGGER_STATUS_INTERVAL_CNT	=	CLK_FREQ_KHZ*TRIGGER_STATUS_INTERVAL;

	//  -------------------------------------------------------------------------------------
	//	ref reg & wire
	//  -------------------------------------------------------------------------------------
	reg		[2:0]								trigger_start_shift			= 3'b0;
	wire										trigger_start_rise			;
	reg		[2:0]								pll_lock_shift				= 3'b0;
	wire										pll_lock_rise				;
	reg											enable						= 1'b0;
	reg		[6:0]								trigger_mode_shfit			= 7'b0;
	reg											lval_dly					= 1'b0;
	reg											fval_dly					= 1'b0;
	wire										fval_rise					;
	wire										fval_fall					;
	reg											image_enable_dly			= 1'b0;
	wire										image_enable_fall			;


	reg											trigger_mode_lock			= 1'b0;

	wire										counter_reset				;//��������λ�ź�
	wire	[31:0]								counter_q					;//���������
	wire										trigger_status_reset		;//trigger_status��λ�ź�

	reg											trigger_status				= 1'b0;
	reg											pll_lock_for_trig			= 1'b0;//restart֮�󣬽⴮PLL���ȶ�����
	reg											pll_lock_for_continue		= 1'b0;//restart֮�󣬽⴮PLL���ȶ�����
	reg											image_enable				= 1'b0;//ͼ�����ʹ�ܣ�1-���ͼ��0-�����ͼ��

	reg		[SENSOR_DAT_WIDTH*CHANNEL_NUM-1:0]	pix_data_dly				= 'b0;
	reg		[SENSOR_DAT_WIDTH*CHANNEL_NUM-1:0]	pix_data_reg				= 'b0;
	reg											fval_reg					= 1'b0;
	reg											lval_reg					= 1'b0;


	//	ref ARCHITECTURE

	//  ===============================================================================================
	//	ref create edge
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	i_trigger_start ȡ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		trigger_start_shift	<=	{trigger_start_shift[1:0],i_trigger_start};
	end
	assign		trigger_start_rise	= (trigger_start_shift[2:1]==2'b01);

	//  -------------------------------------------------------------------------------------
	//	i_pll_lock ȡ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		pll_lock_shift	<=	{pll_lock_shift[1:0],i_pll_lock};
	end
	assign		pll_lock_rise	= (pll_lock_shift[2:1]==2'b01);

	//	-------------------------------------------------------------------------------------
	//	ʹ���ź�
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		enable	<= i_acquisition_start & i_stream_enable;
	end

	//  -------------------------------------------------------------------------------------
	//	�г��ź�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_dly	<=	i_fval;
		lval_dly	<=	i_lval;
	end
	assign	fval_rise	= (fval_dly==1'b0 && i_fval==1'b1) ? 1'b1 : 1'b0;
	assign	fval_fall	= (fval_dly==1'b1 && i_fval==1'b0) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//	image_enable
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		image_enable_dly	<= image_enable;
	end
	assign	image_enable_fall	= {image_enable_dly,image_enable}==2'b10;

	//  ===============================================================================================
	//	ref trigger mode
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	trigger_mode ��ʱ
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		trigger_mode_shfit	<=	{trigger_mode_shfit[5:0],i_trigger_mode};
	end
	//  -------------------------------------------------------------------------------------
	//	trigger_mode_lock
	//	�ڳ������ڼ�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(i_fval==1'b0 && trigger_status==1'b0) begin
			trigger_mode_lock	<= trigger_mode_shfit[6];
		end
	end

	//  -------------------------------------------------------------------------------------
	//	������ƣ���ֹtrigger_status=1ʱ����ʧ�����ģ���쳣
	//	�ӷ�������DSPʱ��32bit�ӷ�
	//	-------------------------------------------------------------------------------------
	binary_counter binary_counter_inst (
	.clk				(clk					),
	.sclr				(counter_reset			),
	.q					(counter_q				)
	);

	//�� trigger_status Ϊ0 ���� ��������ʱ�򣬼ӷ�������
	assign	counter_reset			= (trigger_status==1'b0 || (counter_q==TRIGGER_STATUS_INTERVAL_CNT)) ? 1'b1 : 1'b0;
	//������������ʱ�� trigger_status ��λ
	assign	trigger_status_reset	= (counter_q==TRIGGER_STATUS_INTERVAL_CNT) ? 1'b1 : 1'b0;

	//  ===============================================================================================
	//	ref cut one frame in trigger mode
	//  ===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	trigger_status �ߵ�ƽ������ʱ���ʾ �Ӵ����źŷ��� �� һ֡ͼ�������
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		//	-------------------------------------------------------------------------------------
		//	trigger_status=1����1100ms����trigger_status��0
		//	-------------------------------------------------------------------------------------
		if(trigger_status_reset) begin
			trigger_status	<=	1'b0;
		end
		//	-------------------------------------------------------------------------------------
		//	i2c��ʼ���ͣ���trigger_status������Ϊ1����ʾ�߼����봥��״̬
		//	-------------------------------------------------------------------------------------
		else if(trigger_start_rise) begin
			trigger_status	<=	1'b1;
		end
		//	-------------------------------------------------------------------------------------
		//	�ڳ������ڼ���ͣ�ɵ�ʱ����trigger_status��0���жϴ�������
		//	���ع�ʱ���£������ź�֮�����ع�ʱ��ͣ�ɣ���Ҫ����ֹͣ
		//	-------------------------------------------------------------------------------------
		else if(i_fval==1'b0 && enable==1'b0) begin
			trigger_status	<=	1'b0;
		end
		//	-------------------------------------------------------------------------------------
		//	����֡�����Ϻ�trigger_status��Ϊ0
		//	-------------------------------------------------------------------------------------
		else if(image_enable_fall) begin
			trigger_status	<=	1'b0;
		end
	end

	//	-------------------------------------------------------------------------------------
	//	pll_lock_for_trig
	//	i2c restart����ͺ󣬽⴮PLL��lock���ͣ���ʱ���ǽ�PLL��λ1ms����λ����������ȶ�������״̬��
	//	ͨ�������trigger_status=1ʱ���⴮PLL��lock�źų��������أ�����Ϊ�⴮PLL�ȶ�������
	//	���ź�ֻ�ڴ���״̬����Ч
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(trigger_status) begin
			if(pll_lock_rise) begin
				pll_lock_for_trig		<=	1'b1;
			end
		end
		else begin
			pll_lock_for_trig		<=	1'b0;
		end
	end

	//	-------------------------------------------------------------------------------------
	//	pll_lock_for_continue
	//	���ź���Ϊ�˽������������ʱ��֡������
	//	������������ʱ�򣬻ᷢ�� restart sensor �����PLL��ʧ����
	//	���������ģʽ�£�Ҫ���� pll lock rise ������Ϊ��һ������֡
	//	����ģʽ�¿���Ҳ����restart�Ĳ������̼���һ�׿��ɵ����̣�ͨ���̼������������˲�֡
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!trigger_mode_lock) begin
			if(pll_lock_rise) begin
				pll_lock_for_continue		<=	1'b1;
			end
		end
		else begin
			pll_lock_for_continue		<=	1'b0;
		end
	end

	//	-------------------------------------------------------------------------------------
	//	image_enable ͼ��ʹ���ź�
	//	����ģʽ�£�һֱΪ1
	//	����ģʽ�£�ץȡ�����ź�֮��ĵ�һ������֡
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		//	-------------------------------------------------------------------------------------
		//	����ģʽ�£�ֻҪpll lock�й�һ�������أ���һֱΪ��
		//	-------------------------------------------------------------------------------------
		if(!trigger_mode_lock) begin
			if(pll_lock_for_continue) begin
				image_enable	<=	1'b1;
			end
			else begin
				image_enable	<=	1'b0;
			end
		end
		//	-------------------------------------------------------------------------------------
		//	����ģʽ�£�Ҫץȡsensor restart ֮��ĵ�һ������֡
		//	1.pll_lock_for_trig==1 ��ʾ�����ź��Ѿ���������pll lock�Ѿ���������
		//	2.fval rise==1 ��ʾpll lock֮����һ������֡���ˣ����������Ҫץȡ�ĵ�һ������֡
		//	3.fval fall==1 ��ʾһ�������Ѿ�����
		//	-------------------------------------------------------------------------------------
		else begin
			if(pll_lock_for_trig) begin
				if(fval_rise) begin
					image_enable	<=	1'b1;
				end
				else if(fval_fall) begin
					image_enable	<=	1'b0;
				end
			end
			else begin
				image_enable	<=	1'b0;
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	ref output
	//  -------------------------------------------------------------------------------------
	//	-------------------------------------------------------------------------------------
	//	��������ź����
	//	-------------------------------------------------------------------------------------
	assign	o_trigger_mode		= trigger_mode_lock;
	assign	o_trigger_status	= trigger_status;

	//  -------------------------------------------------------------------------------------
	//	�������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(i_fval==1'b1 && i_lval==1'b1) begin
			pix_data_dly	<=	iv_pix_data;
		end
	end

	always @ (posedge clk) begin
		if(fval_dly & lval_dly & image_enable) begin
			pix_data_reg	<=	pix_data_dly;
		end
		else begin
			pix_data_reg	<=	{SENSOR_DAT_WIDTH*CHANNEL_NUM{1'b1}};
		end
	end
	assign	ov_pix_data	= pix_data_reg;

	//	-------------------------------------------------------------------------------------
	//	�г��ź����
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_reg	<=	fval_dly & image_enable;
		lval_reg	<=	lval_dly & image_enable;
	end
	assign	o_fval	= fval_reg;
	assign	o_lval	= lval_reg;


endmodule