//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : wrap_frame_buf_traffic
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/6/10 11:03:31	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//`include			"wrap_frame_buf_traffic_def.v"
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module wrap_frame_buf_traffic (
	input			clk		,
	input			reset	,
	input			i_fval	,
	input			i_dval	,
	input	[22:0]	iv_frame_size	,
	output	[31:0]	ov_image_dout	,

	input			i_buf_empty	,
	output			o_buf_rd	,
	input	[32:0]	iv_image_din	,
	output			o_good_frame	,
	output			o_bad_frame
	
);

//	ref signals



//	ref ARCHITECTURE

	//  -------------------------------------------------------------------------------------
	//	���ݲ����߼�
	//  -------------------------------------------------------------------------------------
	wrap_wr_data wrap_wr_data_inst (
	.clk			(clk			),
	.reset			(reset			),
	.i_fval			(i_fval			),
	.i_dval			(i_dval			),
	.iv_frame_size	(iv_frame_size	),
	.ov_image_dout	(ov_image_dout	)
	);

	//  -------------------------------------------------------------------------------------
	//	��֡�������ݵ�ģ��
	//  -------------------------------------------------------------------------------------
	wrap_rd_data wrap_rd_data_inst (
	.clk			(clk		),
	.reset			(reset		),
	.i_buf_empty	(i_buf_empty	),
	.o_buf_rd		(o_buf_rd		),
	.iv_frame_size	(iv_frame_size	),
	.iv_image_din	(iv_image_din	),
	.o_good_frame	(o_good_frame	),
	.o_bad_frame	(o_bad_frame	)
	);



endmodule
