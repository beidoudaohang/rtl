//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : test_image
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/12/4 13:41:28	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ����ͼģ�飬�������ֲ���ͼ
//              1)  : �Ҷ�ֵ����
//						��֡ͼ����һ������ֵ����8bitÿ֡����1��������255ʱ����һ����Ϊ0��
//              2)  : ��̬б����(0-255б����)
//						ÿһ���У����ش����ҵ�������8bitÿ�����ص���1��������255ʱ����һ����Ϊ0��
//						��һ�����ص����ֵ��ȫ0��
//              2)  : ��̬б����(0-255����б����)
//						��0-255б�������ƣ�ֻ��ÿһ֡����ÿ�����ص��������8bitÿ�����ص���1��������255ʱ����һ����Ϊ0��
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module test_image # (
	parameter	SENSOR_DAT_WIDTH	= 10		//sensor ���ݿ��
	)
	(
	//Sensor�����ź�
	input								clk					,	//����ʱ��
	input								i_fval				,	//���ź�
	input								i_lval				,	//���ź�
	input	[SENSOR_DAT_WIDTH-1:0]		iv_pix_data			,	//ͼ������
	//�Ĵ�������
	input	[2:0]						iv_test_image_sel	,	//����ͼѡ��Ĵ���,000:��ʵͼ,001:����ͼ��1�Ҷ�ֵ֡����,110:����ͼ��2��ֹ��б����,010:����ͼ��3������б����
	//���
	output								o_fval				,	//����Ч��o_fval��o_lval����λҪ��֤���������λһ��
	output								o_lval				,	//����Ч
	output	[SENSOR_DAT_WIDTH-1:0]		ov_pix_data				//ͼ������
	);

	//	ref signals
	reg									fval_dly			= 1'b0;
	wire								fval_fall			;
	reg									lval_dly			= 1'b0;
	wire								lval_fall			;
	reg		[7:0]						frame_cnt			= 8'b0;
	reg		[7:0]						line_cnt			= 8'b0;
	reg		[7:0]						col_cnt				= 8'b0;
	reg		[SENSOR_DAT_WIDTH-1:0]		pix_data_reg		= {SENSOR_DAT_WIDTH{1'b0}};

	//	ref ARCHITECTURE


	//  ===============================================================================================
	//	ref ***��ȡ����***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	fval ��ȡ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_dly	<= i_fval;
	end
	assign	fval_fall	= (fval_dly==1'b1 && i_fval==1'b0) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//	lval ��ȡ����
	//	1.�����볡�ź���Чʱ���������ź�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(i_fval) begin
			lval_dly	<= i_lval;
		end
		else begin
			lval_dly	<= 1'b0;
		end
	end
	assign	lval_fall	= (lval_dly==1'b1 && i_lval==1'b0) ? 1'b1 : 1'b0;

	//  ===============================================================================================
	//	ref ***��Ҫ����������***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	֡������
	//	1.������ͼ�Ĵ���=000ʱ����ʵͼ��frame_cnt��λΪȫ0��
	//	2.������ͼ�Ĵ���=001ʱ���Ҷ�ֵ��������ͼ��frame_cnt��λΪȫ0��
	//	3.������ͼ�Ĵ���=110ʱ��0-255��̬б���Ʋ���ͼ��frame_cnt��λΪȫ0��
	//	4.������ͼ�Ĵ���=010ʱ��0-255����б���Ʋ���ͼ����i_fval�½��ص�ʱ��frame_cnt����1��

	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		case(iv_test_image_sel)
			3'b000,3'b001,3'b110	: frame_cnt	<= 2'b00;
			3'b010	: begin
				if(fval_fall) begin
					frame_cnt	<= frame_cnt + 1'b1;
				end
			end
			default	: frame_cnt	<= 2'b00;
		endcase
	end

	//  -------------------------------------------------------------------------------------
	//	�м�����
	//	1.������ͼ�Ĵ���=000ʱ����ʵͼ��line_cnt=frame_cnt��
	//	2.������ͼ�Ĵ���=001ʱ���Ҷ�ֵ��������ͼ��line_cnt=frame_cnt��
	//	3.������ͼ�Ĵ���=110ʱ��0-255��̬б���Ʋ���ͼ����i_fval=0ʱ��line_cnt=frame_cnt����i_fval=1ʱ����i_lval���½��ص���1��
	//	4.������ͼ�Ĵ���=010ʱ��0-255����б���Ʋ���ͼ����i_fval=0ʱ��line_cnt=frame_cnt����i_fval=1ʱ����i_lval���½��ص���1��

	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		case(iv_test_image_sel)
			3'b000,3'b001	: line_cnt	<= frame_cnt;
			3'b110,3'b010	: begin
				if(!i_fval) begin
					line_cnt	<= frame_cnt;
				end
				else begin
					if(lval_fall) begin
						line_cnt	<= line_cnt + 1'b1;
					end
				end
			end
			default		: line_cnt	<= frame_cnt;
		endcase
	end

	//  -------------------------------------------------------------------------------------
	//	�м�����
	//	1.������ͼ�Ĵ���=000ʱ����ʵͼ��col_cnt=line_cnt��
	//	2.������ͼ�Ĵ���=001ʱ���Ҷ�ֵ��������ͼ��i_fval�½���ʱcol_cnt����1��
	//	3.������ͼ�Ĵ���=110ʱ��0-255��̬б���Ʋ���ͼ��i_fval=1ʱ��i_lval=1ʱ��col_cnt����1����������£�col_cnt=line_cnt��
	//	4.������ͼ�Ĵ���=010ʱ��0-255����б���Ʋ���ͼ��i_fval=1ʱ��i_lval=1ʱ��col_cnt����1����������£�col_cnt=line_cnt��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		case(iv_test_image_sel)
			3'b000	: col_cnt	<= line_cnt;
			3'b001	: begin
				if(fval_fall) begin
					col_cnt	<= col_cnt + 1'b1;
				end
			end
			3'b110,3'b010	: begin
				if(i_fval&i_lval) begin
					col_cnt	<= col_cnt + 1'b1;
				end
				else begin
					col_cnt	<= line_cnt;
				end
			end
			default		: col_cnt	<= line_cnt;
		endcase
	end

	//  ===============================================================================================
	//	ref ***���***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	ѡ���������
	//	1.��������г��źŶ���Чʱ
	//	--1.1�������ʵͼ�����������=��������
	//	--1.2����ǲ���ͼ������������еĸ�8bit�ò������ݴ��棬��λ���0������Ľ�βģ�飬��ѵ�λ��ȡ���������Ҫ���ڸ�λ
	//	2.��������г��ź���һ����Чʱ����������Ϊ0
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(i_fval==1'b1 && i_lval==1'b1) begin
			if(iv_test_image_sel==3'b000) begin
				pix_data_reg	<= iv_pix_data;
			end
			else begin
				pix_data_reg	<= {col_cnt[7:0],{(SENSOR_DAT_WIDTH-8){1'b0}}};
			end
		end
		else begin
			pix_data_reg	<= {SENSOR_DAT_WIDTH{1'b0}};
		end
	end

	//  -------------------------------------------------------------------------------------
	//	������ݣ��г��źţ���ʱ����1��
	//  -------------------------------------------------------------------------------------
	assign	ov_pix_data			= pix_data_reg;
	assign	o_fval				= fval_dly;
	assign	o_lval				= lval_dly;



endmodule
