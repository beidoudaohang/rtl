//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : fval_lval_phase
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/4/10 14:13:37	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module fval_lval_phase # (
	parameter			DATA_WIDTH	= 8			//���ݿ��
	)
	(
	input						clk			,	//ʱ��
	input						reset		,	//��λ
	input						i_fval		,	//����Ч
	input						i_lval		,	//����Ч
	input	[DATA_WIDTH-1:0]	iv_din		,	//��������
	output						o_fval		,	//����Ч
	output						o_lval		,	//����Ч
	output	[DATA_WIDTH-1:0]	ov_dout			//�������
	);

	//	ref signals
	reg		[5:0]					fval_shift		= 6'b0;
	reg		[2:0]					lval_shift		= 3'b0;
	reg		[DATA_WIDTH-1:0]		pix_data_dly0	= {DATA_WIDTH{1'b0}};
	reg		[DATA_WIDTH-1:0]		pix_data_dly1	= {DATA_WIDTH{1'b0}};
	reg		[DATA_WIDTH-1:0]		pix_data_dly2	= {DATA_WIDTH{1'b0}};
	
	
	//	ref ARCHITECTURE

	//  -------------------------------------------------------------------------------------
	//	�����г��źź����ݣ�ʹ֮����
	//  -------------------------------------------------------------------------------------
	//	-------------------------------------------------------------------------------------
	//	���ź��ܹ���ʱ6��
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_shift	<= {fval_shift[4:0],i_fval};
	end

	//	-------------------------------------------------------------------------------------
	//	���ź��ܹ���ʱ3��
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		lval_shift	<= {lval_shift[1:0],i_lval};
	end

	//	-------------------------------------------------------------------------------------
	//	�����ź��ܹ���ʱ3��
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		pix_data_dly0	<= iv_din;
		pix_data_dly1	<= pix_data_dly0;
		pix_data_dly2	<= pix_data_dly1;
	end

	assign	o_fval		= fval_shift[5] & i_fval;
	assign	o_lval		= lval_shift[2];
	assign	ov_dout		= pix_data_dly2;



endmodule
