//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : fifo_ctrl
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2013/6/13 10:17:01	:|  ��ʼ�汾
//  -- �Ϻ���       :| 2015/3/30 15:39:19	:|  ������Ľ���module��fifo_con��Ϊfifo_ctrl
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :	ǰ��FIFO�ĸ�λģ�飬����1CLK�ĸ�λ�ź�
//              1)  : �첽FIFO�Ķ�д�˿���Ҫ�Ը�λ�ź�ͬ����������ڸ���ʱ�����3�������ڣ�FIFO���ǳ��ڸ�λ״̬
//
//              2)  : fval��dval֮��Ҫ���㹻�Ŀ�϶
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module fifo_ctrl # (
	parameter		DATA_WIDTH			= 32			//���ݿ��
	(
	input							clk					,	//ʱ������
	input							i_fval				,	//���ź�
	input							i_sval				,	//������Ч�źţ�section_valid
	input	[DATA_WIDTH-1:0]		iv_image_din		,	//ͼ������
	output	[35:0]					ov_front_buf_din	,	//fifoд������
	output							o_reset_front_buf		//ǰ��FIFO��λ�ź�
	);

	//ref signals
	reg				fval_dly		= 1'b0;
	wire			fval_rise		;
	reg				reset_buf_reg	= 1'b0;


	//ref ARCHITECTURE

	//	-------------------------------------------------------------------------------------
	//	��fval�����ص���ʱ����λǰ��FIFO
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_dly		<= i_fval;
	end
	assign	fval_rise	= (fval_dly==1'b0 && i_fval==1'b1) ? 1'b1 : 1'b0;

	//	-------------------------------------------------------------------------------------
	//	svalȡ����
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		sval_dly		<= i_sval;
	end
	assign	sval_rise	= (sval_dly==1'b0 && i_sval==1'b1) ? 1'b1 : 1'b0;

	//	-------------------------------------------------------------------------------------
	//	�������źŴ�һ�ģ���Ϊbuf�ĸ�λ�ź�
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		reset_buf_reg	<= fval_rise;
	end
	assign	o_reset_front_buf	= reset_buf_reg;


endmodule
