//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : pulser_filter_wr
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/2/11 14:43:36	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : дramģ��
//              1)  : ѭ��д4��ram
//
//              2)  : ���뵱ǰ���ڴ�����У���Ҫ��rdģ����������ݶ���
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module pulser_filter_wr # (
	parameter					SENSOR_DAT_WIDTH	= 10		//sensor ���ݿ��
	)
	(
	input								clk					,	//����ʱ��
	input								i_fval				,	//���źţ�i_fval���±�����i_lval���10��ʱ������
	input								i_lval				,	//���ź�
	input	[SENSOR_DAT_WIDTH-1:0]		iv_pix_data			,	//ͼ������
	output	[3:0]						ov_buffer_wr_en		,	//ramдʹ��
	output	[11:0]						ov_buffer_wr_addr	,	//ramд��ַ
	output	[9:0]						ov_buffer_wr_din	,	//ramд����
	output	[SENSOR_DAT_WIDTH-1:0]		ov_lower_line			//��ǰ��������ݣ���������֮����rdģ�������2�����ݶ���
	);

	//	ref signals
	reg									lval_dly			= 1'b0;
	wire								lval_fall			;
	reg		[1:0]						lval_cnt			= 2'b0;
	reg		[3:0]						buffer_wr_en		= 4'b0;
	reg		[11:0]						buffer_wr_addr		= 12'b0;
	reg		[SENSOR_DAT_WIDTH-1:0]		buffer_wr_din_dly0	= {SENSOR_DAT_WIDTH{1'b0}};
	reg		[SENSOR_DAT_WIDTH-1:0]		buffer_wr_din_dly1	= {SENSOR_DAT_WIDTH{1'b0}};
	reg		[SENSOR_DAT_WIDTH-1:0]		buffer_wr_din_dly2	= {SENSOR_DAT_WIDTH{1'b0}};


	//	ref ARCHITECTURE

	//	===============================================================================================
	//	ref ***ȡ����***
	//	===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	�ж�lval�ı���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		lval_dly	<= i_lval;
	end
	assign	lval_fall	= (lval_dly==1'b1 && i_lval==1'b0) ? 1'b1 : 1'b0;

	//	===============================================================================================
	//	ref ***ѭ��дram***
	//	===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	lval���ؼ�����
	//	1.��������ʱ������������
	//	2.������Ч�ǣ�ÿ��һ�У�����������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!i_fval) begin
			lval_cnt	<= 2'b00;
		end
		else begin
			if(lval_fall) begin
				lval_cnt	<= lval_cnt + 1'b1;
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	bufferд�ź�
	//	1.��֡����ʱ��дʹ������
	//	2.��֡��Чʱ�������кţ�ѭ��д��4��ram�С���һ��д��ram0
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!i_fval) begin
			buffer_wr_en	<= 4'b0000;
		end
		else begin
			case(lval_cnt)
				2'b00	: buffer_wr_en	<= {3'b000,i_lval};
				2'b01	: buffer_wr_en	<= {2'b00,i_lval,1'b0};
				2'b10	: buffer_wr_en	<= {1'b0,i_lval,2'b00};
				2'b11	: buffer_wr_en	<= {i_lval,3'b000};
				default	: buffer_wr_en	<= 4'b0000;
			endcase
		end
	end
	assign	ov_buffer_wr_en	= buffer_wr_en;

	//  -------------------------------------------------------------------------------------
	//	bufferд��ַ
	//	1.ÿ�н�����д��ַ����
	//	2.д��ַ ���� lval_dly��������ΪҪ�ͺ�дʹ��1��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!lval_dly) begin
			buffer_wr_addr	<= 12'h0;
		end
		else begin
			buffer_wr_addr	<= buffer_wr_addr + 1'b1;
		end
	end
	assign	ov_buffer_wr_addr	= buffer_wr_addr;

	//  -------------------------------------------------------------------------------------
	//	bufferд����
	//	1.i_lval����һ����Ϊдʹ�ܣ�����ҲҪ��Ӧ�Ĵ�һ��
	//	2.û���õ�������λ����λ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		buffer_wr_din_dly0	<= iv_pix_data;
	end
	assign	ov_buffer_wr_din	= {{(10-SENSOR_DAT_WIDTH){1'b0}},buffer_wr_din_dly0};

	//	===============================================================================================
	//	ref ***�����ǰд����***
	//	===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	�����ӳ�֮���bufferд���ݣ�Ŀ������rdģ����������ݶ���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		buffer_wr_din_dly1	<= buffer_wr_din_dly0;
		buffer_wr_din_dly2	<= buffer_wr_din_dly1;
	end
	assign	ov_lower_line	= buffer_wr_din_dly2;



endmodule
