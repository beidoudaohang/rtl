//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : mt9p031_if
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/10/20 15:44:47	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : �� mer-500-14u3x sync buffer�е���mt9p031�ӿ���صĲ�����ȡ���������ھ���ʱ�ӡ�ʹ�ܺ�����
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module mt9p031_if # (
	parameter	SENSOR_DAT_WIDTH	= 10		//sensor ���ݿ��
	)
	(
	//Sensorʱ����
	input								clk_sensor_pix		,	//sensor���������ʱ��,72Mhz,�뱾��72MhzͬƵ����ͬ�࣬����Ϊ��ȫ�첽�������źţ����sensor��λ��sensorʱ�ӿ���ֹͣ��������ڲ�ʱ�Ӳ�ֹͣ
	input								i_fval				,	//sensor����ĳ���Ч�źţ���clk_sensor_pix�����ض��룬i_fval��������i_lval�½��ض��룬i_fval�½�������i_lval�½��ض���
	input								i_lval				,	//sensor���������Ч�źţ���clk_sensor_pix�����ض��룬i_fval��������i_lval�½��ض��룬i_fval�½�������i_lval�½��ض��룬i_fval��Ч�ڼ�Ҳ�п������
	input	[SENSOR_DAT_WIDTH-1:0]		iv_pix_data			,	//sensor�����ͼ�����ݣ���clk_sensor_pix�����ض��룬��·����10��������
	//����ź�
	input								o_clk_sensor_pix	,	//��������Ч
	output								o_fval				,	//����Ч������Ч
	output								o_lval				,	//����Ч������Ч
	output	[SENSOR_DAT_WIDTH-1:0]		ov_pix_data				//ͼ������
	);

	//	ref signals
	//	-------------------------------------------------------------------------------------
	//	���ز���
	//	1.Sensor��������Ĭ�ϲ�ʹ��idelay���ڣ���Ϊ�ⲿ��·��ʱ�Ѿ����úܺ�
	//	2.Sensor��������idelay ��ֵĬ��Ϊ0
	//	3.��ʱ����ת����FIFO������ѡ��BRAM����DRAM�����18�����16��
	//	-------------------------------------------------------------------------------------
	localparam			SENSOR_DAT_IDELAY_EN		= 0		;	//idelayʹ��
	localparam			SENSOR_DAT_IDELAY_VALUE		= 0		;	//idelay��ʱֵ

	wire	[SENSOR_DAT_WIDTH-1:0]			wv_pix_data_delay	;
	wire									w_fval_delay	;
	wire									w_lval_delay	;
	wire									clk_sensor_pix_bufg	;
	wire									clk_sensor_pix_bufg_inv	;

	reg		[SENSOR_DAT_WIDTH-1:0]			pix_data_iob	= 'b0;
	reg										fval_iob		= 1'b0;
	reg										lval_iob		= 1'b0;

	//	ref ARCHITECTURE
	//  ===============================================================================================
	//	ref ***����Sensor����***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	�����ʱ�� ���� ͬ���ź� ��idelay��ʱ ѡ���Ա����ģ��
	//  -------------------------------------------------------------------------------------
	idelay_top # (
	.SENSOR_DAT_WIDTH			(SENSOR_DAT_WIDTH			),
	.SENSOR_DAT_IDELAY_EN		(SENSOR_DAT_IDELAY_EN		),
	.SENSOR_DAT_IDELAY_VALUE	(SENSOR_DAT_IDELAY_VALUE	)
	)
	idelay_top_inst (
	.iv_pix_data				(iv_pix_data		),
	.i_fval						(i_fval				),
	.i_lval						(i_lval				),
	.ov_pix_data_delay			(wv_pix_data_delay	),
	.o_fval_delay				(w_fval_delay		),
	.o_lval_delay				(w_lval_delay		)
	);

	//  -------------------------------------------------------------------------------------
	//	��·ʱ����ȫ��ʱ����Դ���壬ȫ�ֻ�����֮�������������Է���ʱ���������źŵ�skew
	//  -------------------------------------------------------------------------------------
	BUFG bufg_inst (
	.I	(clk_sensor_pix			),
	.O	(clk_sensor_pix_bufg	)
	);
	assign	clk_sensor_pix_bufg_inv	= !clk_sensor_pix_bufg;

	//  -------------------------------------------------------------------------------------
	//	��IOB��ʹ��register���������԰���ʱ���������������λ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk_sensor_pix_bufg_inv) begin
		pix_data_iob	<= wv_pix_data_delay;
		fval_iob		<= w_fval_delay;
		lval_iob		<= w_lval_delay;
	end

	//	-------------------------------------------------------------------------------------
	//	���
	//	-------------------------------------------------------------------------------------
	assign	o_clk_sensor_pix	= clk_sensor_pix_bufg_inv;
	assign	o_fval				= fval_iob;
	assign	o_lval				= lval_iob;
	assign	ov_pix_data			= pix_data_iob;


	//	-------------------------------------------------------------------------------------
	//	����Ϊ UCF ʾ��Լ������Ҫ�ֶ���ӵ� UCF �У��� RTL �����в���Ҫ��������Ϊ��ʾ
	//	-------------------------------------------------------------------------------------
	//	##	-------------------------------------------------------------------------------------
	//	##	-- ref clk constraint
	//	##	-------------------------------------------------------------------------------------
	//	NET "clk_sensor_pix" TNM_NET = "TNM_clk_sensor_pix";
	//	TIMESPEC "TS_clk_sensor_pix" = PERIOD "TNM_clk_sensor_pix" 72 MHz HIGH 50 %;
	//
	//	##	-------------------------------------------------------------------------------------
	//	##	-- ref input constraint
	//	##	-------------------------------------------------------------------------------------
	//	##	-------------------------------------------------------------------------------------
	//	##	sensor����ӿ�Լ��
	//	##	sensor����Ƶ����72MHz��UI��������13.8ns���Ӳ��Բ���������ǰ����������4.5ns
	//	##	-------------------------------------------------------------------------------------
	//	INST "iv_pix_data<?>"	TNM = "TNM_IN_SENSOR";
	//	INST "i_fval"			TNM = "TNM_IN_SENSOR";
	//	INST "i_lval"			TNM = "TNM_IN_SENSOR";
	//	TIMEGRP "TNM_IN_SENSOR" OFFSET = IN 4 ns VALID 8 ns BEFORE "clk_sensor_pix" FALLING;
	//
	//
	//	INST "data_channel_inst/sync_buffer_inst/pix_data_iob_*" 	IOB=TRUE;
	//	INST "data_channel_inst/sync_buffer_inst/fval_iob" 			IOB=TRUE;
	//	INST "data_channel_inst/sync_buffer_inst/lval_iob" 			IOB=TRUE;

endmodule
