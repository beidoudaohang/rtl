//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : ad_clock_unit
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/8/9 13:15:39	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module ad_clock_unit # (
	parameter	CLK_UNIT_VENDOR		= "xilinx"		//����ʱ��������"xilinx" "lattice"
	)
	(
	input			cli			,
	output			clk			,
	output			clk_ser		,
	output			reset_ser
	);

	//	ref signals
	wire			cli_delay	;
	wire			lock	;

	//	ref ARCHITECTURE

	//	-------------------------------------------------------------------------------------
	//	tCLIDLY typ value is 5 ns
	//	-------------------------------------------------------------------------------------
	assign	#5 cli_delay		= cli;

	//	-------------------------------------------------------------------------------------
	//	����ʱ��
	//	-------------------------------------------------------------------------------------
	generate
		if(CLK_UNIT_VENDOR=="xilinx") begin
			dcm_ad dcm_ad_inst (
			.clk_in		(cli_delay		),
			.dcm_reset	(1'b0			),
			.clk0_out	(clk			),
			.clk_fx_out	(clk_ser		),
			.locked		(lock			)
			);
			assign	reset_ser	= !lock;
		end
		else if(CLK_UNIT_VENDOR=="lattice") begin
			pll_ad pll_ad_inst (
			.CLKI	(cli	),
			.CLKOP	(clk_ser	),
			.CLKOS	(clk		),
			.LOCK	(lock		)
			);
			assign	reset_ser	= !lock;
		end
	endgenerate



endmodule
