//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : wrap_wr_logic
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2013/6/14 14:00:40	:|  ��ʼ�汾
//  -- ��ǿ         :| 2014/11/27 10:16:54	:|  ��ֲ��MER-U3V���̣����ݲ�ƷҪ���ʵ��޸�
//  -- ��ǿ         :| 2015/10/15 17:22:35	:|  ��port����չΪ64bit���
//  -- �Ϻ���       :| 2016/9/14 16:25:07	:|  ��ROI�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :	֡����ģ�鶥��
//						1�����֡ͼ��ǰ��FIFO����д��Ͷ�����MCBP2������д��Ĺ���
//						2�����дָ�루ͼ���������ַ�任��д��ַ���ֽڼ������任�Լ�����������������
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------
module wrap_wr_logic # (
	parameter	DATA_WD										= 64		,	//�������λ������ʹ��ͬһ���
	parameter	DDR3_MEM_DENSITY							= "1Gb"		,	//DDR3 ���� "2Gb" "1Gb" "512Mb"
	parameter	DDR3_MASK_SIZE								= 8			,	//mask size
	parameter	BURST_SIZE									= 32		,	//BURST_SIZE��С
	parameter	WR_FLAG_NUM									= 5			,	//дflag�ĸ���
	parameter	PTR_WIDTH									= 2			,	//��дָ���λ��1-���1֡ 2-���3֡ 3-���7֡ 4-���15֡ 5-���31֡ ... 16-���65535֡
	parameter	BYTE_ADDR_WIDTH								= 27		,	//��Ч��ַλ��DDR3������ͬ��λ��ͬ
	parameter	WR_ADDR_WIDTH   							= 19		,	//֡�ڵ�ַλ��
	parameter	WORD_CNT_WIDTH								= 5			,	//word cnt λ��
	parameter	MCB_BURST_BYTE_NUM_WIDTH					= 8			,	//MCB BYTE ADDR ��λΪ0�ĸ���
	parameter	SENSOR_MAX_WIDTH							= 1280		,	//Sensor��������Ч���
	parameter	LEADER_START_ADDR							= 0			,	//leader���׵�ַ
	parameter	TRAILER_START_ADDR							= 2			,	//trailer���׵�ַ
	parameter	CHUNK_START_ADDR							= 4			,	//chunk���׵�ַ
	parameter	IMAGE_START_ADDR							= 6			,	//image���׵�ַ
	parameter	TRAILER_FINAL_START_ADDR					= 254		,	//trailer_final���׵�ַ
	parameter	REG_WD  						 			= 32			//�Ĵ���λ��
	)
	(
	//	===============================================================================================
	//	ͼ������ʱ����
	//	===============================================================================================
	//  -------------------------------------------------------------------------------------
	//  ͼ����������
	//  -------------------------------------------------------------------------------------
	input							clk_in								,	//ǰ��FIFOд������ʱ��
	input							i_fval								,	//����Ч�źţ�����Ч��clk_inʱ����,i_fval��������Ҫ��i_dval����������ǰ��i_fval���½���Ҫ��i_dval���½����ͺ�i_fval��i_dval������֮��Ҫ���㹻�Ŀ�϶����Сֵ��MAX(6*clk_in,6*clk_frame_buf)��i_fval��i_dval�½���֮��Ҫ���㹻�Ŀ�϶����Сֵ��1*clk_in + 7*clk_frame_buf
	input							i_dval								,	//������Ч�źţ�����Ч��clk_inʱ����������Ч�������ź�һ�������������Ƕ������ź�
	input							i_leader_flag						,	//ͷ����־
	input							i_trailer_flag						,	//β����־
	input							i_chunk_flag						,	//chunk��־
	input							i_image_flag						,	//ͼ���־
	input							i_trailer_final_flag				,	//���һ��trailer
	input	[DATA_WD-1:0]			iv_din								,	//ͼ�����ݣ�64λ��clk_inʱ����
	output							o_front_fifo_overflow				,	//֡��ǰ��FIFO��� 0:֡��ǰ��FIFOû����� 1:֡��ǰ��FIFO���ֹ����������
	//	===============================================================================================
	//	֡���湤��ʱ����
	//	===============================================================================================
	//  -------------------------------------------------------------------------------------
	//  �� wrap_rd_logic ����
	//  -------------------------------------------------------------------------------------
	input							clk									,	//MCB
	input							reset								,	//��λ�ź�
	output	[PTR_WIDTH-1:0]			ov_wr_ptr							,	//дָ��,��֡Ϊ��λ
	output	[WR_ADDR_WIDTH-1:0]		ov_wr_addr							,	//P2������ʹ���źţ���־д��ַ�Ѿ���Ч�����ٲñ�֤�£������ܹ�д��DDR�����źŶԵ�ַ�жϷǳ���Ҫ
	output							o_wr_ptr_changing					,	//дָ�����ڱ仯�źţ��������ģ�飬��ʱ��ָ�벻�ܱ仯
	input	[PTR_WIDTH-1 :0]		iv_rd_ptr							,	//��ָ��,��֡Ϊ��λ
	input							i_reading							,	//���ڶ���־
	output							o_writing							,	//����д��־
	input							i_chunk_mode_active					,	//������Чʱ������
	//  -------------------------------------------------------------------------------------
	//  ��������
	//  -------------------------------------------------------------------------------------
	input							i_stream_enable						,	//��ֹͣ�źţ�clkʱ�����ź���Чʱ������������֡д��֡�棬��Чʱ����ֹͣд�룬����λ��д��ַָ�룬��֡��
	input	[PTR_WIDTH-1:0]			iv_frame_depth						,	//֡������� ������Ϊ 1 - 31.
	output	[PTR_WIDTH-1:0]			ov_frame_depth						,	//֡������� ������Ϊ 1 - 31.������Чʱ���ġ�
	//  -------------------------------------------------------------------------------------
	//  MCB�˿�
	//  -------------------------------------------------------------------------------------
	input							i_calib_done						,	//MCBУ׼����źţ�����Ч��ʱ����δ֪
	output							o_wr_cmd_en							,	//MCB CMD FIFO д�źţ�����Ч
	output	[2:0]					ov_wr_cmd_instr						,	//MCB CMD FIFO ָ��
	output	[5:0]					ov_wr_cmd_bl						,	//MCB CMD FIFO ͻ������
	output	[29:0]					ov_wr_cmd_byte_addr					,	//MCB CMD FIFO ��ʼ��ַ
	input							i_wr_cmd_empty						,	//MCB CMD FIFO ���źţ�����Ч
	input							i_wr_cmd_full						,	//MCB CMD FIFO ���źţ�����Ч
	output							o_wr_en								,	//MCB WR FIFO д�źţ�����Ч
	output	[DDR3_MASK_SIZE-1:0]	ov_wr_mask							,	//MCB WR �����ź�
	output	[DATA_WD-1:0]			ov_wr_data							,	//MCB WR FIFO д����
	input							i_wr_full								//MCB WR FIFO ���źţ�����Ч
	);



	//	ref signals

	localparam	MAX_LINE_DATA				= SENSOR_MAX_WIDTH*2;			//BIT10 12 ģʽ�� һ�е�������
	localparam	MIN_FRONT_FIFO_DEPTH		= MAX_LINE_DATA/(DATA_WD/8);	//ǰ��fifo��ȵ���Сֵ
	localparam	FRONT_FIFO_DEPTH			= (MIN_FRONT_FIFO_DEPTH<=256) ? 256 : ((MIN_FRONT_FIFO_DEPTH<=512) ? 512 : ((MIN_FRONT_FIFO_DEPTH<=1024) ? 1024 : 2048));
	localparam	WR_FLAG_WIDTH				= log2(WR_FLAG_NUM);

	//FSM Parameter Define
	parameter	S_IDLE		= 3'd0;
	parameter	S_PTR		= 3'd1;
	parameter	S_WR		= 3'd2;
	parameter	S_CMD		= 3'd3;
	parameter	S_FLAG		= 3'd4;

	reg		[2:0]	current_state	= S_IDLE;
	reg		[2:0]	next_state		= S_IDLE;

	//FSM for sim
	// synthesis translate_off
	reg		[127:0]			state_ascii;
	always @ ( * ) begin
		case(current_state)
			3'd0 :	state_ascii	<= "S_IDLE";
			3'd1 :	state_ascii	<= "S_PTR";
			3'd2 :	state_ascii	<= "S_WR";
			3'd3 :	state_ascii	<= "S_CMD";
			3'd4 :	state_ascii	<= "S_FLAG";
		endcase
	end
	// synthesis translate_on

	//	-------------------------------------------------------------------------------------
	//	ȡ��������ȡ��
	//	-------------------------------------------------------------------------------------
	function integer log2 (input integer xx);
		integer x;
		begin
			x	= xx-1 ;
			for (log2=0;x>0;log2=log2+1) begin
				x	= x >> 1;
			end
		end
	endfunction

	//	-------------------------------------------------------------------------------------
	//	��̬λ��ƴ��
	//	1.����verilog�е�λ��ƴ��������в�������ֱ����������function�ķ�ʽʵ�ֶ�̬λ��ƴ��
	//	-------------------------------------------------------------------------------------
	//	i		              ptr_and_addr
	//
	//	i=0		        |------------------------|
	//	i=1		        ||-----------------------|
	//	i=2		        | |----------------------|
	//	i=3		        |  |---------------------|
	//	i=4		        |   |--------------------|
	//	i=5		        |    |-------------------|
	//                    ^           ^
	//			        |ptr |       addr        |
	//	-------------------------------------------------------------------------------------
	//	for ѭ��չ��֮��
	//  -------------------------------------------------------------------------------------
	//	i		���֡��	frame_depth��Χ		byte_addrʵ���Ų�
	//	i=0		1			1					{{(30-WR_ADDR_WIDTH-MCB_BURST_BYTE_NUM_WIDTH){1'b0}},wr_addr[WR_ADDR_WIDTH-1:0],{(MCB_BURST_BYTE_NUM_WIDTH){1'b0}}}
	//	i=1		2			2       			{{(30-WR_ADDR_WIDTH-MCB_BURST_BYTE_NUM_WIDTH){1'b0}},wr_ptr[0:0],wr_addr[WR_ADDR_WIDTH-2:0],{(MCB_BURST_BYTE_NUM_WIDTH){1'b0}}}
	//	i=2		4			3-4					{{(30-WR_ADDR_WIDTH-MCB_BURST_BYTE_NUM_WIDTH){1'b0}},wr_ptr[1:0],wr_addr[WR_ADDR_WIDTH-3:0],{(MCB_BURST_BYTE_NUM_WIDTH){1'b0}}}
	//	i=3 	8			5-8					{{(30-WR_ADDR_WIDTH-MCB_BURST_BYTE_NUM_WIDTH){1'b0}},wr_ptr[2:0],wr_addr[WR_ADDR_WIDTH-4:0],{(MCB_BURST_BYTE_NUM_WIDTH){1'b0}}}
	//	i=4		16			9-16				{{(30-WR_ADDR_WIDTH-MCB_BURST_BYTE_NUM_WIDTH){1'b0}},wr_ptr[3:0],wr_addr[WR_ADDR_WIDTH-5:0],{(MCB_BURST_BYTE_NUM_WIDTH){1'b0}}}
	//	i=5		32			17-32				{{(30-WR_ADDR_WIDTH-MCB_BURST_BYTE_NUM_WIDTH){1'b0}},wr_ptr[4:0],wr_addr[WR_ADDR_WIDTH-6:0],{(MCB_BURST_BYTE_NUM_WIDTH){1'b0}}}
	//	i=6		64			33-64				{{(30-WR_ADDR_WIDTH-MCB_BURST_BYTE_NUM_WIDTH){1'b0}},wr_ptr[5:0],wr_addr[WR_ADDR_WIDTH-7:0],{(MCB_BURST_BYTE_NUM_WIDTH){1'b0}}}
	//	i=7		128			65-128				{{(30-WR_ADDR_WIDTH-MCB_BURST_BYTE_NUM_WIDTH){1'b0}},wr_ptr[6:0],wr_addr[WR_ADDR_WIDTH-8:0],{(MCB_BURST_BYTE_NUM_WIDTH){1'b0}}}
	//	i=8		256			129-256				{{(30-WR_ADDR_WIDTH-MCB_BURST_BYTE_NUM_WIDTH){1'b0}},wr_ptr[7:0],wr_addr[WR_ADDR_WIDTH-9:0],{(MCB_BURST_BYTE_NUM_WIDTH){1'b0}}}
	//	......
	//	-------------------------------------------------------------------------------------
	function [WR_ADDR_WIDTH-1:0] ptr_and_addr;
		input	[PTR_WIDTH-1:0]	ptr_int;
		input	[WR_ADDR_WIDTH-1:0]	addr_int;
		input	[PTR_WIDTH-1:0]	depth_int;
		integer	i;
		integer	j;
		begin
			if(depth_int==1) begin
				ptr_and_addr	= addr_int;
			end
			for(i=1;i<=PTR_WIDTH;i=i+1) begin
				if(depth_int>=(2**(i-1)+1) && depth_int<=2**i) begin
					for(j=0;j<WR_ADDR_WIDTH;j=j+1) begin
						if(j<WR_ADDR_WIDTH-i) begin
							ptr_and_addr[j]	= addr_int[j];
						end
						else begin
							ptr_and_addr[j]	= ptr_int[j+i-WR_ADDR_WIDTH];
						end
					end
				end
			end
		end
	endfunction



	reg		[2:0]						fval_shift			= 3'b000;
	wire								fval_rise			;
	wire								fval_fall			;
	reg									stream_enable_reg	= 1'b0;
	reg		[1:0]						calib_done_shift	= 2'b00;
	reg									active_flag_dly		= 1'b0;
	wire								active_flag_fall	;
	reg		[PTR_WIDTH-1:0]				frame_depth_reg 	= 'b0;
	wire								reset_fifo			;
	wire								fifo_wr_en			;
	wire								fifo_full			;
	wire	[DATA_WD+4:0]				fifo_din			;
	wire								fifo_rd_en			;
	reg									front_fifo_overflow	= 1'b0;
	reg									wr_cmd_en			= 1'b0;
	wire	[WR_ADDR_WIDTH-1:0]			ptr_and_addr_int	;
	wire								fifo_empty			;
	wire								fifo_prog_empty		;
	wire	[DATA_WD+4:0]				fifo_dout			;

	reg		[PTR_WIDTH-1:0]				wr_ptr				= 'b0;
	reg		[WR_ADDR_WIDTH-1:0]			wr_addr				= 'b0;
	reg		[WORD_CNT_WIDTH-1:0]		word_cnt 			= {(WORD_CNT_WIDTH){1'b1}};
	reg									able_to_write 		= 1'b0;
	wire								leader_flag			;
	wire								trailer_flag		;
	wire								chunk_flag			;
	wire								image_flag			;
	wire								trailer_final_flag	;
	wire								active_flag			;
	reg		[WR_FLAG_WIDTH-1:0]			flag_num_cnt		= 'b0;
	wire	[BYTE_ADDR_WIDTH-1:0]		start_addr			;
	reg									wr_ptr_changing		= 1'b0;
	reg									writing_reg			= 1'b0;



	//	ref ARCHITECTURE


	//	===============================================================================================
	//	ref ***edge***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	fval ������
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_shift	<= {fval_shift[1:0],i_fval};
	end
	assign	fval_rise	= (fval_shift[2:1]==2'b01) ? 1'b1 : 1'b0;
	assign	fval_fall	= (fval_shift[2:1]==2'b10) ? 1'b1 : 1'b0;

	//	-------------------------------------------------------------------------------------
	//	stream_enable_reg
	//	1.�� i_stream_enable =0ʱ��������Ϊ0
	//	2.�� i_stream_enable =1 �� fval rise ��ʱ�򣬲��ܱ�Ϊ1
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(i_stream_enable==1'b0) begin
			stream_enable_reg	<= 1'b0;
		end
		else if(fval_rise==1'b1) begin
			stream_enable_reg	<= 1'b1;
		end
	end

	//	-------------------------------------------------------------------------------------
	//	i_calib_done ʱ����δ֪����Ҫ��2�Ĵ���
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		calib_done_shift	<= {calib_done_shift[0],i_calib_done};
	end

	//	-------------------------------------------------------------------------------------
	//	��ǰѡ�е�flag�ı���
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		active_flag_dly	<= active_flag;
	end
	assign	active_flag_fall	= (active_flag_dly==1'b1 && active_flag==1'b0) ? 1'b1 : 1'b0;

	//	-------------------------------------------------------------------------------------
	//	frame_depth_reg ֡����ȼĴ���
	//	1.�ڿ���״̬���� frame_depth
	//	2.�����0���򱣻�Ϊ1
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(current_state==S_IDLE) begin
			if(iv_frame_depth==0) begin
				frame_depth_reg	<= 1;
			end
			else begin
				frame_depth_reg	<= iv_frame_depth;
			end
		end
	end
	assign	ov_frame_depth	= frame_depth_reg;

	//	===============================================================================================
	//	ref ***front fifo***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	front fifo ����
	//	-------------------------------------------------------------------------------------
	generate
		//	-------------------------------------------------------------------------------------
		//	sensor�п�С�ڵ���1024
		//	-------------------------------------------------------------------------------------
		if(FRONT_FIFO_DEPTH==256) begin
			frame_buf_front_fifo_w69d256_pe128 frame_buf_front_fifo_w69d256_pe128_inst (
			.rst			(reset_fifo			),
			.wr_clk			(clk_in				),
			.wr_en			(fifo_wr_en			),
			.full			(fifo_full			),
			.din			(fifo_din			),
			.rd_clk			(clk				),
			.rd_en			(fifo_rd_en			),
			.empty			(fifo_empty			),
			.prog_empty		(fifo_prog_empty	),
			.dout			(fifo_dout			)
			);
		end
		//	-------------------------------------------------------------------------------------
		//	sensor�п�С�ڵ���2048
		//	-------------------------------------------------------------------------------------
		else if(FRONT_FIFO_DEPTH==512) begin
			frame_buf_front_fifo_w69d512_pe256 frame_buf_front_fifo_w69d512_pe256_inst (
			.rst			(reset_fifo			),
			.wr_clk			(clk_in				),
			.wr_en			(fifo_wr_en			),
			.full			(fifo_full			),
			.din			(fifo_din			),
			.rd_clk			(clk				),
			.rd_en			(fifo_rd_en			),
			.empty			(fifo_empty			),
			.prog_empty		(fifo_prog_empty	),
			.dout			(fifo_dout			)
			);
		end
		//	-------------------------------------------------------------------------------------
		//	sensor�п�С�ڵ���4096
		//	-------------------------------------------------------------------------------------
		else if(FRONT_FIFO_DEPTH==1024) begin
			frame_buf_front_fifo_w69d1024_pe512 frame_buf_front_fifo_w69d1024_pe512_inst (
			.rst			(reset_fifo			),
			.wr_clk			(clk_in				),
			.wr_en			(fifo_wr_en			),
			.full			(fifo_full			),
			.din			(fifo_din			),
			.rd_clk			(clk				),
			.rd_en			(fifo_rd_en			),
			.empty			(fifo_empty			),
			.prog_empty		(fifo_prog_empty	),
			.dout			(fifo_dout			)
			);
		end
		//	-------------------------------------------------------------------------------------
		//	sensor�п�С�ڵ���8192
		//	-------------------------------------------------------------------------------------
		else if(FRONT_FIFO_DEPTH==2048) begin
			frame_buf_front_fifo_w69d2048_pe1024 frame_buf_front_fifo_w69d2048_pe1024_inst (
			.rst			(reset_fifo			),
			.wr_clk			(clk_in				),
			.wr_en			(fifo_wr_en			),
			.full			(fifo_full			),
			.din			(fifo_din			),
			.rd_clk			(clk				),
			.rd_en			(fifo_rd_en			),
			.empty			(fifo_empty			),
			.prog_empty		(fifo_prog_empty	),
			.dout			(fifo_dout			)
			);
		end
	endgenerate

	//	-------------------------------------------------------------------------------------
	//	fifo ��λ
	//	1.ʱ�Ӹ�λ fval������ ͣ��ֱ��fval������ ������������ÿһ�����ܹ���λ
	//	2.�첽fifo�ĸ�λ�źſ���������ʱ����ģ���Ϊ��fifo�ڲ�������ͬ�������˴����źŶ���clkʱ����ġ�
	//	-------------------------------------------------------------------------------------
	assign	reset_fifo	= reset | fval_rise | !stream_enable_reg;

	//	-------------------------------------------------------------------------------------
	//	fifo дʹ��
	//	clk_inʱ�����ڳ��źš������ź���Ч��ʱ����fifo������ʱ�򣬲���д
	//	-------------------------------------------------------------------------------------
	assign	fifo_wr_en	= i_fval & i_dval & !fifo_full;

	//	-------------------------------------------------------------------------------------
	//	fifo ��������
	//	1.fifo�������ݹ���69bit����5bit��flag����64bit������
	//	-------------------------------------------------------------------------------------
	assign	fifo_din	= {i_trailer_final_flag,i_image_flag,i_chunk_flag,i_trailer_flag,i_leader_flag,iv_din};

	//  -------------------------------------------------------------------------------------
	//  FIFO ���ź�
	//	1.������д״̬ʱ�����ǰ��fifo���գ���fifo�����������ź���Ч����ǰflag��Ч������ź���Ч
	//	2.������߼�����������ᵼ�¶��������
	//  -------------------------------------------------------------------------------------
	assign	fifo_rd_en	= (current_state==S_WR) & !fifo_empty & !i_wr_full & stream_enable_reg & active_flag;

	//	-------------------------------------------------------------------------------------
	//	֡��ǰ��������
	//	1.һ������ǰ��fifo��������������Ϊ1��û�а취��λ�����������ϵ�
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk_in) begin
		if(fifo_wr_en && fifo_full) begin
			front_fifo_overflow <= 1'b1;
		end
	end
	assign o_front_fifo_overflow = front_fifo_overflow;

	//	===============================================================================================
	//	ref ***mcb fifo operation***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	mcb wr fifo дʹ���ź���fifo�Ķ�ʹ���ź���ͬһ��
	//	-------------------------------------------------------------------------------------
	assign	o_wr_en		= fifo_rd_en;

	//	-------------------------------------------------------------------------------------
	//	û��mask��byte��ȫ��Ҫд�뵽fifo��
	//	-------------------------------------------------------------------------------------
	assign	ov_wr_mask	= 'b0;

	//	-------------------------------------------------------------------------------------
	//	дָ��
	//	1.���ݲ������壬������2�����ʽ
	//	2.3'b010 -> with precharge; 3'b000 -> without precharge
	//	-------------------------------------------------------------------------------------
	assign	ov_wr_cmd_instr	= 3'b000;

	//	-------------------------------------------------------------------------------------
	//	MCB CMD FIFO д�ź�
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		//	-------------------------------------------------------------------------------------
		//	������ CMD ״̬ʱ�����cmd fifo�������Ϳ���д��һ���µ�����
		//	-------------------------------------------------------------------------------------
		if((current_state==S_CMD && i_wr_cmd_full==1'b0)) begin
			wr_cmd_en	<= 1'b1;
		end
		//	-------------------------------------------------------------------------------------
		//	������ FLAG ״̬ʱ�����cmd fifo�������Ϳ���д��һ���µ�����
		//	-------------------------------------------------------------------------------------
		else if(current_state==S_FLAG && i_wr_cmd_full==1'b0 && wr_cmd_en==1'b0) begin
			wr_cmd_en	<= 1'b1;
		end
		else begin
			wr_cmd_en	<= 1'b0;
		end
	end
	assign	o_wr_cmd_en	= wr_cmd_en;

	//  -------------------------------------------------------------------------------------
	//  MCB fifo д����
	//	1.ǰ��FIFO���ֱ���͵�MCB��fifo��
	//	2.ǰ��FIFO���� first word fall through���ص㣬�����յ�ʱ�򣬵�һ�������Ѿ��ŵ��˿�����
	//	3.��ǰ��FIFO��MCB WR FIFO֮��û�м���ˮ�ߣ�Ŀ���Ǽ�����Դ��ʵ�������ﲢ�����ǹؼ�·��������Ҫ���ġ�
	//  -------------------------------------------------------------------------------------
	assign	ov_wr_data	= fifo_dout[DATA_WD-1:0];

	//	-------------------------------------------------------------------------------------
	//	д����
	//	1.burst_length=word_cnt����ͼ���ва���ʱ�򣬲��Ὣ���������д��DDR
	//	2.��ͣ�ɵ�ʱ��д��64�����ݣ�Ŀ���Ǳ�֤���п�ͣ�ɲ����������� mcb wr fifo
	//	-------------------------------------------------------------------------------------
	assign	ov_wr_cmd_bl	= (stream_enable_reg==1'b1) ? {{(6-WORD_CNT_WIDTH){1'b0}},word_cnt} : 6'b111111;

	//  -------------------------------------------------------------------------------------
	//	mcb ��ַƴ��
	//	1.UG388 pg63 �Ե�ַ�ֲ�����ϸ������
	//	2.burst_size ��С��ͬ�����λ�̶�Ϊ0�ĸ���Ҳ��ͬ
	//	3.���� iv_frame_depth ����˿�λ����16������֧�ֵ���󻺴����Ϊ2**16-1=65535֡
	//	4.���ݵ�ǰ�趨��֡������ȣ����ı�洢λ��
	//	-------------------------------------------------------------------------------------
	assign	ptr_and_addr_int	= ptr_and_addr(wr_ptr[PTR_WIDTH-1:0],wr_addr[WR_ADDR_WIDTH-1:0],frame_depth_reg[PTR_WIDTH-1:0]);
	assign	ov_wr_cmd_byte_addr	= {{(30-WR_ADDR_WIDTH-MCB_BURST_BYTE_NUM_WIDTH){1'b0}},ptr_and_addr_int[WR_ADDR_WIDTH-1:0],{(MCB_BURST_BYTE_NUM_WIDTH){1'b0}}};

	//	===============================================================================================
	//	ref ***ptr addr cnt***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	дָ���߼�
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		//	-------------------------------------------------------------------------------------
		//	��֡�������1֡���߸�λ�ź���Ч����ʹ����Чʱ��дָ�븴λ
		//	-------------------------------------------------------------------------------------
		if(frame_depth_reg==1 || reset==1'b1 || stream_enable_reg==1'b0) begin
			wr_ptr	<= 0;
		end
		else begin
			//	-------------------------------------------------------------------------------------
			//	ֻ���� PTR ״̬�� wr_ptr_changing=1��ʱ�򣬲��ܸı�дָ��
			//	-------------------------------------------------------------------------------------
			if(current_state==S_PTR && wr_ptr_changing==1'b1) begin
				//	-------------------------------------------------------------------------------------
				//	�����ڶ���ʱ��дָ�벻�ܽ����ָ��
				//	-------------------------------------------------------------------------------------
				if(i_reading==1'b1) begin
					//	-------------------------------------------------------------------------------------
					//	��дָ���Ѿ��ﵽ���ֵʱ
					//	1.�����ģ�����ڶ�0���ڴ棬��ôдָ��Ҫ������ָ�룬ʵ��д��Խ
					//	2.�����ģ��û���ڶ�0���ڴ棬��ôдָ��д0�ŵ�ַ
					//	-------------------------------------------------------------------------------------
					if(wr_ptr==(frame_depth_reg-1)) begin
						if(iv_rd_ptr==0) begin
							wr_ptr	<= 1;
						end
						else begin
							wr_ptr	<= 0;
						end
					end
					//	-------------------------------------------------------------------------------------
					//	��дָ��û�дﵽ���ֵ�����Ƕ�ָ�뵽�����ֵʱ
					//	1.���дָ��+1=��ָ�룬��ôдָ��д0�ŵ�ַ
					//	2.���дָ��+1!=��ָ�룬��ôдָ������
					//	-------------------------------------------------------------------------------------
					else if(iv_rd_ptr==(frame_depth_reg-1)) begin
						if((wr_ptr+1'b1)==iv_rd_ptr) begin
							wr_ptr	<= 0;
						end
						else begin
							wr_ptr	<= wr_ptr + 1'b1;
						end
					end
					//	-------------------------------------------------------------------------------------
					//	�����������дָ�붼�������ֵ
					//	1.���дָ��+1=��ָ�룬��ôдָ��Ҫ������ָ�룬ʵ��д��Խ
					//	2.���дָ��+1!=��ָ�룬��ôдָ������
					//	-------------------------------------------------------------------------------------
					else begin
						if((wr_ptr+1'b1)==iv_rd_ptr) begin
							wr_ptr	<= iv_rd_ptr + 1'b1;
						end
						else begin
							wr_ptr	<= wr_ptr + 1'b1;
						end
					end
				end
				//	-------------------------------------------------------------------------------------
				//	�����ڶ�=0ʱ��˵����ģ��û��ռ���κ��ڴ棬дָ������������
				//	1.���дָ��ﵽ�����ֵ����д0���ڴ�
				//	2.���дָ��û�дﵽ�����ֵ����дָ������
				//	-------------------------------------------------------------------------------------
				else begin
					if(wr_ptr==(frame_depth_reg-1)) begin
						wr_ptr	<= 0;
					end
					else begin
						wr_ptr	<= wr_ptr + 1'b1;
					end
				end
			end
		end
	end
	assign	ov_wr_ptr		= wr_ptr;

	//  -------------------------------------------------------------------------------------
	//  д��ַ�߼�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		//	-------------------------------------------------------------------------------------
		//	��idle״̬�£���ַ����
		//	-------------------------------------------------------------------------------------
		if(current_state==S_IDLE) begin
			wr_addr	<= 'b0;
		end
		//	-------------------------------------------------------------------------------------
		//	��flag״̬�£���д�����֮��д��ַ�л�Ϊ��һ��flag�ĵ�ַ
		//	-------------------------------------------------------------------------------------
		else if(current_state==S_FLAG && wr_cmd_en==1'b1) begin
			wr_addr	<= start_addr[BYTE_ADDR_WIDTH-1:MCB_BURST_BYTE_NUM_WIDTH];
		end
		//	-------------------------------------------------------------------------------------
		//	������״̬�£���д�����֮��д��ַ����
		//	-------------------------------------------------------------------------------------
		else if(wr_cmd_en==1'b1) begin
			wr_addr	<= wr_addr + 1'b1;
		end
	end
	assign	ov_wr_addr	= wr_addr;

	//	-------------------------------------------------------------------------------------
	//	word_cnt һ��burst������
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		//	-------------------------------------------------------------------------------------
		//	1.һ��burst�ļ����������� burst_size
		//	2.����Ҫ���ж�reset����Ϊreset=1���ͻ����idle״̬
		//	3.��һ֡��ʼ��ʱ����ռ���������wr_addrһͬ���㡣
		//	-------------------------------------------------------------------------------------
		if(current_state==S_IDLE) begin
			word_cnt	<= {(WORD_CNT_WIDTH){1'b1}};
		end
		//	-------------------------------------------------------------------------------------
		//	1.��flag״̬��д������Ч����������λ
		//	2.��Ϊ�л�flag��ʱ���п��ܴ�ʱ��word_cnt��û�дﵽ���ֵ�������Ҫ�ֶ�����
		//	-------------------------------------------------------------------------------------
		else if(current_state==S_FLAG && wr_cmd_en==1'b1) begin
			word_cnt	<= {(WORD_CNT_WIDTH){1'b1}};
		end
		//	-------------------------------------------------------------------------------------
		//	��CMD״̬�£��������һ֡�����ˣ���ôҪ��word cnt��λ����wr״̬���ж��Ƿ��idle
		//	-------------------------------------------------------------------------------------
		else if(current_state==S_CMD && fifo_empty==1'b1 && fval_shift[1]==1'b0) begin
			word_cnt	<= {(WORD_CNT_WIDTH){1'b1}};
		end
		//	-------------------------------------------------------------------------------------
		//	���������£�ÿ��һ��ǰ��fifo��word_cnt����
		//	-------------------------------------------------------------------------------------
		else if(fifo_rd_en==1'b1) begin
			word_cnt	<= word_cnt + 1'b1;
		end
	end

	//	-------------------------------------------------------------------------------------
	//	flag ������
	//	-------------------------------------------------------------------------------------
	assign	leader_flag				= fifo_dout[DATA_WD];
	assign	trailer_flag			= fifo_dout[DATA_WD+1];
	assign	chunk_flag				= fifo_dout[DATA_WD+2];
	assign	image_flag				= fifo_dout[DATA_WD+3];
	assign	trailer_final_flag		= fifo_dout[DATA_WD+4];

	//	-------------------------------------------------------------------------------------
	//	active_flag ��ǰѡ�е�flag
	//	-------------------------------------------------------------------------------------
	assign	active_flag		= fifo_dout[DATA_WD+flag_num_cnt];

	//	-------------------------------------------------------------------------------------
	//	flag_num_cnt
	//	��ǰflag�½��ص�ʱ�򣬼���������
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(current_state==S_IDLE) begin
			flag_num_cnt	<= 'b0;
		end
		else if(active_flag_fall) begin
			//	-------------------------------------------------------------------------------------
			//	���chunkû�� ������chunk
			//	-------------------------------------------------------------------------------------
			if(i_chunk_mode_active==1'b0 && flag_num_cnt==1) begin
				flag_num_cnt	<= 3;
			end
			else begin
				flag_num_cnt	<= flag_num_cnt + 1'b1;
			end

		end
	end

	//	-------------------------------------------------------------------------------------
	//	start_addr ÿ��flag����ʼ��ַ ��byteΪ��λ
	//	1.����flag_cnt �жϵ�ǰ������һ��״̬
	//	2.�˴�����ʹ������߼���Ҳ����ʹ��ʱ���߼�������ʵ�ʲ��ߵ����������˴�Ϊ�ؼ�·�������Ը�Ϊʱ���߼���
	//	-------------------------------------------------------------------------------------
	//				________
	//	active_flag	       |____________________
	//				       ___
	//	af_fall		_______| |__________________
	//                         ___
	//	wr_cmd		___________| |______________
	//
	//	flag_num_cnt|  0     |  1               |
	//
	//	state		|  WR  |C| F |  WR          |
	//
	//	start_addr	|  0     |  1               |
	//
	//	word_cnt	|  0         |  1           |
	//
	//	-------------------------------------------------------------------------------------
	assign	start_addr	=
	(flag_num_cnt==0) ? LEADER_START_ADDR : (
	(flag_num_cnt==1) ? TRAILER_START_ADDR : (
	(flag_num_cnt==2) ? CHUNK_START_ADDR : (
	(flag_num_cnt==3) ? IMAGE_START_ADDR : (
	(flag_num_cnt==4) ? TRAILER_FINAL_START_ADDR : (
	LEADER_START_ADDR
	)))));

	//	===============================================================================================
	//	ref ***wr rd communication***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	��״̬������ PTR ״̬��ʱ��wr_ptr_change����Ϊ1������״̬������Ϊ0
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(current_state==S_PTR) begin
			wr_ptr_changing	<= 1'b1;
		end
		else begin
			wr_ptr_changing	<= 1'b0;
		end
	end
	assign	o_wr_ptr_changing	= wr_ptr_changing;

	//  -------------------------------------------------------------------------------------
	//  ����д
	//	1.������idle״̬ʱ������д�ź�����
	//	2.������ PTR ״̬�� wr_ptr_changing=1��ʱ�򣬲��ܱ�Ϊ1������Ҫ�� wr_ptr һ��ı��ԭ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(current_state==S_IDLE) begin
			writing_reg	<= 1'b0;
		end
		else if(current_state==S_PTR && wr_ptr_changing==1'b1) begin
			//	-------------------------------------------------------------------------------------
			//	1.�ڵ�֡ʱ�����һ֡���ڶ���������д��ʹ��
			//	2.��������һ��������������дʹ��
			//	-------------------------------------------------------------------------------------
			if(frame_depth_reg==1 && i_reading==1'b1) begin
				writing_reg	<= 1'b0;
			end
			else begin
				writing_reg	<= 1'b1;
			end
		end
	end
	assign	o_writing	= writing_reg;

	//	===============================================================================================
	//	ref ***FSM***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	FSM Sequential Logic
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(reset) begin
			current_state	<= S_IDLE;
		end
		else begin
			current_state	<= next_state;
		end
	end

	//	-------------------------------------------------------------------------------------
	//	FSM Conbinatial Logic
	//	-------------------------------------------------------------------------------------
	always @ ( * ) begin
		case(current_state)
			S_IDLE	:
			//	-------------------------------------------------------------------------------------
			//	IDLE -> PTR
			//	1.������Ч 2.У׼��� 3.ǰ��fifo���գ�˵������
			//	-------------------------------------------------------------------------------------
			if(stream_enable_reg==1'b1 && calib_done_shift[1]==1'b1 && fifo_empty==1'b0) begin
				next_state	= S_PTR;
			end
			else begin
				next_state	= S_IDLE;
			end
			S_PTR	:
			//	-------------------------------------------------------------------------------------
			//	PTR״̬����ʱ��2��CLK����PTR�ڼ䷢��wr_ptr_change�źţ�wr_ptr_change�źŵ�������2��ʱ������
			//	������ wr_ptr_changing=1��ʱ�򣬿����ж�״̬��ת
			//	PTR -> IDLE
			//	1.�ڵ�֡ʱ�����һ֡���ڶ�������IDLE״̬
			//	PTR -> WR
			//	1.��������ת��IDLE������������ת��WR״̬
			//	-------------------------------------------------------------------------------------
			if(wr_ptr_changing==1'b1) begin
				if(frame_depth_reg==1 && i_reading==1'b1) begin
					next_state	= S_IDLE;
				end
				else begin
					next_state	= S_WR;
				end
			end
			else begin
				next_state	= S_PTR;
			end
			S_WR	:
			//	-------------------------------------------------------------------------------------
			//	WR -> IDLE
			//	1.ǰ��fifo�� 2.fval=0 3.��һ�η���cmd֮��û�д�ǰ��fifo��ȡ����
			//	-------------------------------------------------------------------------------------
			if((fifo_empty==1'b1 && fval_shift[1]==1'b0 && word_cnt==(BURST_SIZE-1)) || (stream_enable_reg==1'b0 && word_cnt==(BURST_SIZE-1))) begin
				next_state	= S_IDLE;
			end
			//	-------------------------------------------------------------------------------------
			//	WR -> CMD
			//	1.��ǰ��fifo�ж������������� BURST_SIZE-2 �� ���ڶ�ǰ��fifo ��
			//	2.ǰ��fifo�� �� fval=0 �� ��ǰ��fifo�ж�ȡ��һ�������� ��
			//	3.ͣ��
			//	-------------------------------------------------------------------------------------
			else if((word_cnt==(BURST_SIZE-2) && fifo_rd_en==1'b1) || (fifo_empty==1'b1 && fval_shift[1]==1'b0 && word_cnt!=(BURST_SIZE-1)) || stream_enable_reg==1'b0) begin
				next_state	= S_CMD;
			end
			//	-------------------------------------------------------------------------------------
			//	WR -> FLAG
			//	1.��ǰflag�½���
			//	-------------------------------------------------------------------------------------
			else if(active_flag_fall==1'b1) begin
				next_state	= S_FLAG;
			end
			else begin
				next_state	= S_WR;
			end
			S_CMD	:
			//	-------------------------------------------------------------------------------------
			//	CMD -> FLAG
			//	1.��ǰflag�½���
			//	-------------------------------------------------------------------------------------
			if(active_flag_fall==1'b1) begin
				next_state	= S_FLAG;
			end
			//	-------------------------------------------------------------------------------------
			//	CMD -> WR
			//	1.��ǰflagû���½���
			//	2.wr cmd fifoû����
			//	-------------------------------------------------------------------------------------
			else if(i_wr_cmd_full==1'b0) begin
				next_state	= S_WR;
			end
			else begin
				next_state	= S_CMD;
			end
			S_FLAG	:
			//	-------------------------------------------------------------------------------------
			//	���뵽FLAG״̬��word cnt�ܿ��ܲ���31�����Ҫ�ֶ���λ������Ҫ��֤д�źź�cmd�źŲ���ͬʱ��Ч
			//	FLAG�Ŀ������2��ʱ�����ڣ�CMD��FLAG�����һ�����ڲ��������� mcb wr fifo en �� mcb wr cmd �Ͳ���ͬʱ��Ч
			//	-------------------------------------------------------------------------------------
			//	-------------------------------------------------------------------------------------
			//	FLAG -> WR
			//	1.wr cmd en ��Ч �� ��ǰ�������һ��flag
			//	-------------------------------------------------------------------------------------
			if(wr_cmd_en==1'b1) begin
				next_state	= S_WR;
			end
			else begin
				next_state	= S_FLAG;
			end
			default	:
			next_state	= S_IDLE;
		endcase
	end


endmodule