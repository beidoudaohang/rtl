//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : harness
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/3/9 17:18:50	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------
`define		TESTCASE	testcase_1
module harness ();

	//	ref signals
	//	===============================================================================================
	//	--ref parameter
	//	===============================================================================================


	//	===============================================================================================
	//	--ref signal
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	����
	//	-------------------------------------------------------------------------------------
	wire							reset		;
	wire							clk			;
	wire	[7:0]					iv_din		;
	wire							i_wr		;
	wire							i_rd		;

	//	-------------------------------------------------------------------------------------
	//	���
	//	-------------------------------------------------------------------------------------
	wire							o_full_sync			;
	wire							o_half_full_sync	;
	wire							o_empty_sync		;
	wire	[7:0]					ov_dout_sync		;

	wire							o_full_bb			;
	wire							o_half_full_bb		;
	wire							o_data_present_bb	;
	wire	[7:0]					ov_dout_bb			;

	//	-------------------------------------------------------------------------------------
	//	����
	//	-------------------------------------------------------------------------------------



	//	ref ARCHITECTURE

	//	-------------------------------------------------------------------------------------
	//	���������ź�
	//	-------------------------------------------------------------------------------------
	assign	clk						= `TESTCASE.clk	;
	assign	reset					= `TESTCASE.reset	;
	assign	iv_din					= `TESTCASE.iv_din	;
	assign	i_wr					= `TESTCASE.i_wr	;
	assign	i_rd					= `TESTCASE.i_rd	;


	//	-------------------------------------------------------------------------------------
	//	���� dut ģ��
	//	-------------------------------------------------------------------------------------
	sync_fifo_srl_w8d16 sync_fifo_srl_w8d16_inst (
	.reset			(reset			),
	.clk			(clk			),
	.iv_din			(iv_din			),
	.i_wr			(i_wr			),
	.o_full			(o_full_sync		),
	.o_half_full	(o_half_full_sync	),
	.ov_dout		(ov_dout_sync	),
	.i_rd			(i_rd			),
	.o_empty		(o_empty_sync	)
	);

	bbfifo_16x8 bbfifo_16x8_inst (
	.reset			(reset			),
	.clk			(clk			),
	.write			(i_wr			),
	.data_in		(iv_din			),
	.full			(o_full_bb		),
	.half_full		(o_half_full_bb	),
	.read			(i_rd			),
	.data_out		(ov_dout_bb		),
	.data_present	(o_data_present_bb	)
	);



	//generate vcd file
	//initial begin
	//$dumpfile("test.vcd");
	//$dumpvars(1,top_frame_buffer_inst);
	//end

	//for lattice simulation
	//GSR   GSR_INST (.GSR (1'b1)); //< global reset sig>
	//PUR   PUR_INST (.PUR (1'b1)); //<powerup reset sig>



endmodule
