//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : map_python
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/10/14 9:55:41	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ����������Ϊpython�������ʽ
//              1)  : AN66427-D д����python������������з�ʽ
//
//						--even kernel--			--odd kernel--
//				ch0		p0			p1			p7			p6
//
//				ch1		p2			p3			p5			p4
//
//				ch2		p4			p5			p3			p2
//
//				ch3		p6			p7			p1			p0
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module map_python # (
	parameter			DATA_WIDTH			= 8		,	//����λ��
	parameter			CHANNEL_NUM			= 4			//ͨ����
	)
	(
	input										clk							,	//ʱ��
	input										i_fval						,	//����Ч
	input										i_lval						,	//����Ч
	input	[DATA_WIDTH*CHANNEL_NUM-1:0]		iv_pix_data					,	//��������
	output										o_fval						,	//����Ч
	output										o_lval						,	//����Ч
	output	[DATA_WIDTH*CHANNEL_NUM-1:0]		ov_pix_data						//��������
	);


	//	ref signals

	reg		[1:0]								pix_cnt	= 2'b0;
	reg		[1:0]								pix_cnt_dly0	= 2'b0;
	reg		[1:0]								pix_cnt_dly1	= 2'b0;
	reg		[1:0]								pix_cnt_dly2	= 2'b0;
	wire	[DATA_WIDTH-1:0]					wv_data_lane	[CHANNEL_NUM-1:0]	;
	reg		[DATA_WIDTH-1:0]					map_temp0	[CHANNEL_NUM-1:0];
	reg		[DATA_WIDTH-1:0]					map_temp1	[CHANNEL_NUM-1:0];
	wire	[DATA_WIDTH*CHANNEL_NUM-1:0]		map_temp_align0	;
	wire	[DATA_WIDTH*CHANNEL_NUM-1:0]		map_temp_align1	;
	reg		[DATA_WIDTH*CHANNEL_NUM-1:0]		map_latch0	;
	reg		[DATA_WIDTH*CHANNEL_NUM-1:0]		map_latch1	;
	reg		[DATA_WIDTH*CHANNEL_NUM-1:0]		dout_reg	= 'b0;
	reg		[3:0]								fval_shift	= 4'b0;
	reg		[3:0]								lval_shift	= 4'b0;



	//	ref ARCHITECTURE
	//	===============================================================================================
	//	ref ***��������***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	���ؼ�����
	//	--8���������1��kernel��2��kernel���һ��ѭ��
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(i_fval&i_lval) begin
			pix_cnt	<= pix_cnt + 1'b1;
		end
		else begin
			pix_cnt	<= 4'b0;
		end
	end


	always @ (posedge clk) begin
		pix_cnt_dly0	<= pix_cnt;
		pix_cnt_dly1	<= pix_cnt_dly0;
		pix_cnt_dly2	<= pix_cnt_dly1;
	end
	//	-------------------------------------------------------------------------------------
	//	����ͨ��
	//	--ÿ��ͨ����λ���� DATA_WIDTH ��bit
	//	--��ˣ���ߵ�ͨ���ڵ�byte��С�ˣ���͵�ͨ���ڵ�byte��
	//	-------------------------------------------------------------------------------------
	genvar	i;
	generate
		for(i=0;i<CHANNEL_NUM;i=i+1) begin
			assign	wv_data_lane[i]	= iv_pix_data[DATA_WIDTH*(i+1)-1:DATA_WIDTH*i];
		end
	endgenerate

	//-------------------------------------------------------------------------------------------------
	//						***input***
	//-------------------------------------------------------------------------------------------------
	//
	//				ch0		p0			p4			p0			p4
	//
	//				ch1		p1			p5			p1			p5
	//
	//				ch2		p2			p6			p2			p6
	//
	//				ch3		p3			p7			p3			p7
	//
	//-------------------------------------------------------------------------------------------------
	//						***output***
	//-------------------------------------------------------------------------------------------------
	//						--even kernel--			--odd kernel--
	//				ch0		p0			p1			p7			p6
	//
	//				ch1		p2			p3			p5			p4
	//
	//				ch2		p4			p5			p3			p2
	//
	//				ch3		p6			p7			p1			p0
	//
	//-------------------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(i_fval&i_lval) begin
			case(pix_cnt)
				0	: begin
					map_temp0[0]		<= wv_data_lane[0];
					map_temp1[0]		<= wv_data_lane[1];
					map_temp0[1]		<= wv_data_lane[2];
					map_temp1[1]		<= wv_data_lane[3];
				end
				1	: begin
					map_temp0[2]		<= wv_data_lane[0];
					map_temp1[2]		<= wv_data_lane[1];
					map_temp0[3]		<= wv_data_lane[2];
					map_temp1[3]		<= wv_data_lane[3];
				end
				2	: begin
					map_temp1[3]		<= wv_data_lane[0];
					map_temp0[3]		<= wv_data_lane[1];
					map_temp1[2]		<= wv_data_lane[2];
					map_temp0[2]		<= wv_data_lane[3];
				end
				3	: begin
					map_temp1[1]		<= wv_data_lane[0];
					map_temp0[1]		<= wv_data_lane[1];
					map_temp1[0]		<= wv_data_lane[2];
					map_temp0[0]		<= wv_data_lane[3];
				end
			endcase
		end
	end

	//	-------------------------------------------------------------------------------------
	//         		  ___  ___  ___  ___  ___  ___  ___  ___  ___  ___  ___  ___  ___  ___  ___  ___  ___  ___  ___  ___  ___  ___
	//	clk  		__| |__| |__| |__| |__| |__| |__| |__| |__| |__| |__| |__| |__| |__| |__| |__| |__| |__| |__| |__| |__| |__| |__
	//
	//					   ________________________________________________________________________________________________
	//	i_fval		_______|                                                                                              |_________
	//                     _________________________________________              _________________________________________
	//	i_lval		_______|                                       |______________|                                       |_________
	//
	//	pix_cnt		-------< 0 >< 1 >< 2 >< 3 >< 0 >< 1 >< 2 >< 3 >< 0            >< 0 >< 1 >< 2 >< 3 >< 0 >< 1 >< 2 >< 3 >
	//
	//	din			-------<d0 ><d1 ><d2 ><d3 ><d4 ><d5 ><d6 ><d7 >----------------<d0 ><d1 ><d2 ><d3 ><d4 ><d5 ><d6 ><d7 >----------------
	//
	//	map_temp0	-----------------<d01><xxx><d23><xxx><d45><xxx><d67><xxx>----------------<d01><xxx><d23><xxx><d45><xxx><d67><xxx>----------------
	//
	//	map_temp1	-----------------<d01><xxx><d23><xxx><d45><xxx><d67><xxx>----------------<d01><xxx><d23><xxx><d45><xxx><d67><xxx>----------------
	//
	//	map_latch0	----------------------<d01     ><d23     ><d45     ><d67     >----------------<d01     ><d23     ><d45     ><d67     >----------------
	//
	//	map_latch1	----------------------<d01     ><d23     ><d45     ><d67     >----------------<d01     ><d23     ><d45     ><d67     >----------------
	//
	//	pix_cnt_dly2----------------------< 0 >< 1 >< 2 >< 3 >< 0 >< 1 >< 2 >< 3 >< 0            >< 0 >< 1 >< 2 >< 3 >< 0 >< 1 >< 2 >< 3 >
	//
	//	dout		---------------------------<d0 ><d1 ><d2 ><d3 ><d4 ><d5 ><d6 ><d7 >----------------<d0 ><d1 ><d2 ><d3 ><d4 ><d5 ><d6 ><d7 >----------------
	//
	//					                       ________________________________________________________________________________________________
	//	o_fval		___________________________|                                                                                              |_________
	//                                         _________________________________________              _________________________________________
	//	o_lval		___________________________|                                       |______________|                                       |_________
	//
	//
	//	-------------------------------------------------------------------------------------


	//	===============================================================================================
	//	ref ***���***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	����ͨ��
	//	--ÿ��ͨ����λ���� DATA_WIDTH ��bit
	//	--��ˣ���ߵ�ͨ���ڵ�byte��С�ˣ���͵�ͨ���ڵ�byte��
	//	-------------------------------------------------------------------------------------
	genvar	j;
	generate
		for(j=0;j<CHANNEL_NUM;j=j+1) begin
			assign	map_temp_align0[DATA_WIDTH*(j+1)-1:DATA_WIDTH*j]	= map_temp0[j];
			assign	map_temp_align1[DATA_WIDTH*(j+1)-1:DATA_WIDTH*j]	= map_temp1[j];
		end
	endgenerate

	//	-------------------------------------------------------------------------------------
	//	�� pix_cnt[0]==0 ʱ���������е�����
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!pix_cnt[0]) begin
			map_latch0	<= map_temp_align0;
			map_latch1	<= map_temp_align1;
		end
	end

	//	-------------------------------------------------------------------------------------
	//	ѡ�����������
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(pix_cnt_dly2[0]) begin
			dout_reg	<= map_latch0;
		end
		else begin
			dout_reg	<= map_latch1;
		end
	end
	assign	ov_pix_data	= dout_reg;

	//	-------------------------------------------------------------------------------------
	//	������ʱ2�ģ�ʹ��ҲҪ��ʱ2��
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_shift	<= {fval_shift[2:0],i_fval};
	end
	assign	o_fval	= fval_shift[3];

	always @ (posedge clk) begin
		lval_shift	<= {lval_shift[2:0],i_lval};
	end
	assign	o_lval	= lval_shift[3];

endmodule
