//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : fix_reg_list
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/3/6 11:24:55	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : fixʱ����ļĴ����б�
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module fix_reg_list # (
	parameter		SPI_ADDR_LENGTH				= 16	,	//spi ��ַ�ĳ���
	parameter		SHORT_REG_WD				= 16	,	//�̼Ĵ���λ��
	parameter		REG_WD						= 32	,	//�Ĵ���λ��
	parameter		LONG_REG_WD					= 64		//���Ĵ���λ��
	)
	(
	//  ===============================================================================================
	//	�����ź�
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	spiʱ����
	//  -------------------------------------------------------------------------------------
	input								i_rd_en			,	//��ʹ�ܣ�clk_sampleʱ����
	input	[SPI_ADDR_LENGTH-1:0]		iv_addr			,	//��д��ַ��clk_sampleʱ����
	//  -------------------------------------------------------------------------------------
	//	�̶���ƽ
	//  -------------------------------------------------------------------------------------
	output								o_fix_sel		,	//�̶�ʱ����ѡ��
	output	[SHORT_REG_WD-1:0]			ov_fix_rd_data		//������
	);

	//	ref signals

	//  ===============================================================================================
	//	ref �汾��
	//  ===============================================================================================
	localparam	VENDOR_ID		= 16'h4448;
	localparam	PRODUCT_ID		= 16'h0000;
	localparam	FPGA_VERSION_H	= 16'h0102;
	localparam	FPGA_VERSION_L	= 16'h0123;
	localparam	TEST_VERSION	= 16'h1001;

	//  ===============================================================================================
	//	���ƼĴ���
	//  ===============================================================================================
	reg		[SHORT_REG_WD:0]			data_out_reg= {(SHORT_REG_WD+1){1'b0}};

	//	ref ARCHITECTURE

	//  ===============================================================================================
	//	ref ***������***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	-- ref �����̼Ĵ�������
	//	��, data_out_reg ���bit˵���Ƿ�ѡ���˸�ʱ������������Ϊ�Ĵ�������
	//  -------------------------------------------------------------------------------------
	always @ ( * ) begin
		//������ַѡ�е�ʱ��pix sel����Ϊ��Ч
		if(i_rd_en) begin
			case(iv_addr[8:0])
				//  -------------------------------------------------------------------------------------
				//	�汾
				//  -------------------------------------------------------------------------------------
				9'h00	: data_out_reg	<= {1'b1,VENDOR_ID};
				9'h01	: data_out_reg	<= {1'b1,PRODUCT_ID};
				9'h02	: data_out_reg	<= {1'b1,FPGA_VERSION_H};
				9'h03	: data_out_reg	<= {1'b1,FPGA_VERSION_L};
				9'h04	: data_out_reg	<= {1'b1,TEST_VERSION};

				default	: data_out_reg	<= {(SHORT_REG_WD+1){1'b0}};

			endcase
		end
		//����ʹ��ȡ����ʱ��sel���ܸ�λΪ0
		else begin
			data_out_reg	<= {(SHORT_REG_WD+1){1'b0}};
		end
	end
	assign	o_fix_sel		= data_out_reg[SHORT_REG_WD];
	assign	ov_fix_rd_data	= data_out_reg[SHORT_REG_WD-1:0];


endmodule