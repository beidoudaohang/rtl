//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : stream_ctrl
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/12/4 16:54:58	:|  ��ʼ�汾
//  -- �Ϻ���       :| 2015/10/21 9:56:38	:|  �� sync_buffer ģ�����������ƹ���
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ���2��������
//              1)  : �Ĵ�����Чʱ��
//						����ͨ�����õļĴ�������Ҫ�����ģ��������Чʱ�����������fval������ʱ�������Ĵ���
//				2)  : ��ͣ�ɿ��ƣ������������֡���Ƶ�ʹ���ź�
//
//				3)  :
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module stream_ctrl # (
	parameter					SENSOR_DAT_WIDTH	= 10	,	//sensor ���ݿ��
	parameter					CHANNEL_NUM			= 4		,	//��������ͨ������
	parameter					REG_WD				= 32		//�Ĵ���λ��
	)
	(
	//����ʱ����
	input											clk					,	//����ʱ����
	input											i_fval				,	//clk_pixʱ����sync buffer�����fval�ź�
	input											i_lval				,	//clk_pixʱ����sync buffer�����lval�ź�
	input	[SENSOR_DAT_WIDTH*CHANNEL_NUM-1:0]		iv_pix_data			,	//clk_pixʱ����sync buffer�����pix data�ź�
	output											o_fval				,	//����Ч��չ��o_fval��o_fval��ǰ���ذ�סl_fvalԼ10��ʱ��
	output											o_lval				,	//����Ч
	output	[SENSOR_DAT_WIDTH*CHANNEL_NUM-1:0]		ov_pix_data			,	//ͼ������
	//�����ź�
	input											i_acquisition_start	,	//�����źţ�0-ͣ�ɣ�1-����
	input											i_stream_enable		,	//��ʹ���ź�
	input											i_encrypt_state		,	//����ͨ·�����dna ʱ���򣬼���״̬�����ܲ�ͨ���������ͼ��
	//�Ĵ�������
	input	[REG_WD-1:0]							iv_pixel_format		,	//���ظ�ʽ�Ĵ���
	input	[2:0]									iv_test_image_sel	,	//����ͼѡ��Ĵ���,000:��ʵͼ,001:����ͼ��1�Ҷ�ֵ֡����,110:����ͼ��2��ֹ��б����,010:����ͼ��3������б����
	//������Чʱ���ļĴ���
	output											o_full_frame_state	,	//����֡״̬,�üĴ���������֤ͣ��ʱ�������֡,0:ͣ��ʱ���Ѿ�������һ֡����,1:ͣ��ʱ�����ڴ���һ֡����
	output	[REG_WD-1:0]							ov_pixel_format		,	//��sync buffer������Чʱ������
	output	[2:0]									ov_test_image_sel		//��sync buffer������Чʱ������
	);

	//	ref signals
	reg												fval_dly			= 1'b0;
	wire											fval_rise			;
	reg												encrypt_state_dly0	= 1'b0;
	reg												encrypt_state_dly1	= 1'b0;
	reg												enable				= 1'b0;
	reg												fval_reg			= 1'b0;
	reg												lval_reg			= 1'b0;
	reg		[SENSOR_DAT_WIDTH*CHANNEL_NUM-1:0]		pix_data_reg		= 8'b0;
	reg												full_frame_state	= 1'b0;
	reg		[REG_WD-1:0]							pixel_format_reg	= {REG_WD{1'b0}};
	reg		[2:0]									test_image_sel_reg	= 3'b000;

	//	ref ARCHITECTURE
	//  ===============================================================================================
	//	ref ***��ʹ�ܿ���***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	fval ȡ����
	//	1.�첽ʱ�����䣬��Ҫ������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_dly	<= i_fval;
	end
	assign	fval_rise	= (fval_dly==1'b0 && i_fval==1'b1) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//	����״̬ͬ��
	//	1.i_encrypt_state�� osc bufgʱ������źţ����β���ͨ����pixʱ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		encrypt_state_dly0	<= i_encrypt_state;
		encrypt_state_dly1	<= encrypt_state_dly0;
	end

	//  -------------------------------------------------------------------------------------
	//	enable ����֡ʹ�ܿ����ź�
	//	1.�� i_fval �� o_fval ���ǵ͵�ƽʱ������enable�Ĵ�����enable=���������ź������״̬������
	//	2.�� i_fval �� o_fval ������1���ߵ�ƽʱ������enable�Ĵ�������֤����֡
	//	3.i_fval=1 o_fval=0ʱ����һ��ʱ�����ڣ�o_fval=1����ʱ������������֡�жϣ���Ϊ��һ�����ڿ϶������fval
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(i_fval==1'b0 && o_fval==1'b0) begin
			enable	<= i_stream_enable & i_acquisition_start & encrypt_state_dly1;
		end
	end

	//  ===============================================================================================
	//	ref ***�������***
	//  ===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	fval reg
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(enable==1'b0) begin
			fval_reg	<= 1'b0;
		end
		else begin
			fval_reg	<= i_fval;
		end
	end
	assign	o_fval	= fval_reg;

	//	-------------------------------------------------------------------------------------
	//	lval reg
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(enable==1'b0) begin
			lval_reg	<= 1'b0;
		end
		else begin
			lval_reg	<= i_lval;
		end
	end
	assign	o_lval	= lval_reg;

	//	-------------------------------------------------------------------------------------
	//	pix_data_reg
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(enable==1'b0) begin
			pix_data_reg	<= 'b0;
		end
		else begin
			pix_data_reg	<= iv_pix_data;
		end
	end
	assign	ov_pix_data	= pix_data_reg;

	//  ===============================================================================================
	//	ref ***��־���Ĵ�������***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	-- ref ����֡��־
	//	1.�� i_stream_enable=0ʱ����������֡��־
	//	2.�� i_fval_sync=0ʱ����������֡��־
	//	3.�� i_fval_sync=1��i_acquisition_start=0ʱ������֡��λ
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!i_stream_enable || !o_fval) begin
			full_frame_state	<= 1'b0;
		end
		else begin
			if(o_fval==1'b1 && i_acquisition_start==1'b0) begin
				full_frame_state	<= 1'b1;
			end
		end
	end
	assign	o_full_frame_state	= full_frame_state;

	//  -------------------------------------------------------------------------------------
	//	-- ref �Ĵ�����Чʱ������
	//	1.��fval_rise=1����һ֡����ʱ�����¼Ĵ���
	//	2.����ʱ�̣��������ظ�ʽ�Ĵ���
	//	3.��Щ�Ĵ�������������ͨ���в�ֹһ��ģ��ʹ�ã����Ҫ������ͨ������ǰ�˿���
	//  -------------------------------------------------------------------------------------
	//	���ظ�ʽ�Ĵ���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(fval_rise) begin
			pixel_format_reg	<= iv_pixel_format;
		end
	end
	assign	ov_pixel_format		= pixel_format_reg;

	//  -------------------------------------------------------------------------------------
	//	����ͼѡ��Ĵ���
	//	--���д����ǷǷ�ֵ��������һ�εĽ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(fval_rise) begin
			if(iv_test_image_sel==3'b000 || iv_test_image_sel==3'b001 || iv_test_image_sel==3'b110 || iv_test_image_sel==3'b010) begin
				test_image_sel_reg	<= iv_test_image_sel;
			end
		end
	end
	assign	ov_test_image_sel		= test_image_sel_reg;

endmodule