//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : bitslip
//  -- �����       : �ܽ�
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �ܽ�       :| 2015/08/11 13:46:45	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ����HiSPiЭ���ͬ���ֶ���word�߽�
//					 �ڽ��ж������ʱ����lane1Ϊ�ο���lane1���ݶ���������laneҲӦ���Ƕ���ġ������
//					 ʵ��������laneû�ж��룬��˵������lane��ʱ�ӵ���λ��ϵ���ԣ�������ݽ�����λ������
//             		 ��Ϊ����������ͬ���֣�������û�м�⵽ͬ����ʱ��ÿ��1�������ڽ���һ�μ�⡣
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ns
//-------------------------------------------------------------------------------------------------
module bitslip # (
	parameter		SER_FIRST_BIT			= "LSB"				,	//"LSB" or "MSB" , first bit to the receiver
	parameter		END_STYLE				= "LITTLE"			,	//"LITTLE" or "BIG" , "LITTLE" - {CHANNEL3 CHANNE2 CHANNEL1 CHANNEL0}. "BIG" - {CHANNEL0 CHANNEL1 CHANNEL2 CHANNEL3}.
	parameter		SENSOR_DAT_WIDTH		= 12				,	//sensor��������λ��
	parameter		RATIO					= 6					,	//�⴮����
	parameter		CHANNEL_NUM				= 4						//ͨ����
	)
	(
	input												clk						,	//���벢��ʱ��
	input												reset					,	//����ʱ����λ�ź�
	input	[RATIO*CHANNEL_NUM-1:0]						iv_data					,	//���벢������
	input	[15:0]										iv_line_length			,	//������
	input												i_bitslip_en			,	//bitslipʹ�ܣ�Ϊ�ߵ�ƽʱ���ж������
	output												o_bitslip				,	//���bitslipʹ�ܣ�����selectIO
	output												o_data_valid			,	//ͨ��������Ч�ź�
	output												o_clk_en				,	//ʱ��ʹ���ź�
	output	[SENSOR_DAT_WIDTH*CHANNEL_NUM-1:0]			ov_data						//�Ѿ�����������
	);

	//ref signals

	//	-------------------------------------------------------------------------------------
	//	hispi ��ͬ����
	//	--����LSBʱ���Ƚ��յ��Ͱ��ֽڣ������λ�Ĵ��������ơ��������ȳ�����word���������档ͬ������36'h000_000_fff��
	//	--����MSBʱ���Ƚ��յ��Ͱ��ֽڣ������λ�Ĵ��������ơ��������ȳ�����word���������档ͬ������36'hfff_000_000��
	//	-------------------------------------------------------------------------------------
	localparam	SYNC_WORD	= (END_STYLE=="LITTLE") ? {{4*RATIO{1'b0}},{2*RATIO{1'b1}}} : {{2*RATIO{1'b1}},{4*RATIO{1'b0}}};

	reg		[1:0]									bitslip_en_shift		;	//��λʹ�ܴ�����
	wire	[RATIO-1:0]								wv_data_lane[CHANNEL_NUM-1:0]	;	//������ϵ�ͨ��1������
	reg		[2*RATIO-1:0]							data_lane_align[CHANNEL_NUM-1:0]	;	//������ϵ�ͨ��1������
	reg												div_cnt					= 1'b0	;	//��Ƶ������
	reg		[RATIO*6-1:0]							data_lane0_shift		= 'b0	;	//lan0ͨ����λ�Ĵ���

	reg												data_lock				= 'b0	;	//�߽�����־λ��1��ʾ�߽��Ѿ�����
	reg		[15:0]									bitslip_cnt				= 'b0	;	//�����������ÿ�������ڽ���һ�ζ������
	reg												bitslip_reg				= 1'b0	;	//iserdes��λʹ���ź�

	//ref ARCHITECTURE
	//	===============================================================================================
	//	ref ***�첽ʱ������***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	i_bitslip_enΪclk_pixʱ����ת����i_clk_parallelʱ����
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk)begin
		bitslip_en_shift	<=	{bitslip_en_shift[0],i_bitslip_en};
	end

	//	===============================================================================================
	//	ref ***���ͬ����***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	����ͨ��
	//	--ÿ��ͨ����λ���� RATIO ��bit
	//	--��ˣ���ߵ�ͨ���ڵ�byte��С�ˣ���͵�ͨ���ڵ�byte��
	//	-------------------------------------------------------------------------------------
	genvar	i;
	generate
		for(i=0;i<CHANNEL_NUM;i=i+1) begin
			if(END_STYLE=="LITTLE") begin
				assign	wv_data_lane[i]	= iv_data[RATIO*(i+1)-1:RATIO*i];
			end
			else if(END_STYLE=="BIG") begin
				assign	wv_data_lane[i]	= iv_data[RATIO*(CHANNEL_NUM-i)-1:RATIO*(CHANNEL_NUM-i-1)];
			end
		end
	endgenerate

	//	-------------------------------------------------------------------------------------
	//	��lan0��λ��ÿ���ƶ� RATIO ��bit
	//	--Ŀǰ�ļ�ⷽ����ֻ��lane0���ͬ���֡�����ͨ�������
	//	--lan0�� RATIO bit����ÿ����λ��ע�⣬�˴�������LSB MSB �����ǽ����ݴ���Ͷ��Ƶ���߶�
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(SER_FIRST_BIT=="LSB") begin
			data_lane0_shift	<= {wv_data_lane[0],data_lane0_shift[RATIO*6-1:RATIO]};
		end
		else if(SER_FIRST_BIT=="MSB") begin
			data_lane0_shift	<= {data_lane0_shift[RATIO*5-1:0],wv_data_lane[0]};
		end
	end

	//	-------------------------------------------------------------------------------------
	//	���ͬ����
	//	--��⵽{{L{1'b1}},{L{1'b0}},{L{1'b0}}}���ʾ��⵽ͬ���֣�ͬʱ�߽�Ҳ�Ƕ����
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk)begin
		if(reset==1'b1 || bitslip_en_shift[1]==1'b0)begin
			data_lock	<=	0;
		end
		else begin
			if(data_lane0_shift[RATIO*6-1:0]==SYNC_WORD)begin
				data_lock	<=	1;
			end
		end
	end

	//	-------------------------------------------------------------------------------------
	//	��LSBΪ����˵��data lock��ƴ���߼�
	//	-------------------------------------------------------------------------------------
	//	-------------------------------------------------------------------------------------
	//			  	  ____   ____   ____   ____   ____   ____   ____   ____   ____   ____   ____   ____   ____   ____
	//	clk_2x		__|  |___|  |___|  |___|  |___|  |___|  |___|  |___|  |___|  |___|  |___|  |___|  |___|  |___|  |___
	//
	//	byte in		--<L0    ><H0   ><L1   ><H1   ><L2   ><H2   ><L3   ><H3   ><L4   ><H4   ><L5   ><H5   ><L6   ><H6   >
	//
	//									                 ______________________________________________________________________
	//	data lock	_____________________________________|
	//
	//	byte shift	------------------------------<L0H0L1H1>
	//
	//	data align	-------------------------------------<L2H1  ><H2L2 ><L3H2 ><H3L3 ><L4H3 ><H4L4 ><L5H4 ><H5L5 ><L6H5 >
	//						    								________      ________      ________      ________
	//	clk en		____________________________________________|      |______|      |______|      |______|      |______
	//
	//
	//	-------------------------------------------------------------------------------------

	//	===============================================================================================
	//	ref ***ƴ������***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	ÿ��ͨ������ʱ1��
	//	--2�� RATIO bit��ƴ��һ��word
	//	--LSBģʽ���Ƚ��յ��� RATIO bit�ǵ�λ��MSBģʽ���Ƚ��յ��� RATIO bit�Ǹ�λ
	//	-------------------------------------------------------------------------------------
	genvar	j;
	generate
		for(j=0;j<CHANNEL_NUM;j=j+1) begin
			if(SER_FIRST_BIT=="LSB") begin
				always @ (posedge clk) begin
					data_lane_align[j]	= {wv_data_lane[j],data_lane_align[j][2*RATIO-1:RATIO]};
				end
			end
			else if(SER_FIRST_BIT=="MSB") begin
				always @ (posedge clk) begin
					data_lane_align[j]	= {data_lane_align[j][RATIO-1:0],wv_data_lane[j]};
				end
			end
		end
	endgenerate

	//	-------------------------------------------------------------------------------------
	//	div_cnt ��Ƶ������
	//	--ֻ�� data_lock == 1��ʱ��ſ�ʼ����
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!data_lock) begin
			div_cnt	<= 'b0;
		end
		else begin
			div_cnt	<= !div_cnt;
		end
	end
	assign	o_clk_en	= div_cnt;

	//	===============================================================================================
	//	ref ***bitslip ����߼�***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	�����ڼ�����
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk)begin
		if(reset==1'b1 || bitslip_en_shift[1]==1'b0)begin
			bitslip_cnt	<=	'd0;
		end
		else begin
			if(bitslip_cnt==iv_line_length) begin
				bitslip_cnt	<= 'b0;
			end
			else begin
				bitslip_cnt	<= bitslip_cnt + 1'b1;
			end
		end
	end

	//	-------------------------------------------------------------------------------------
	//	��һ��֮��û�м�⵽ͬ���֣�����λ
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(reset==1'b1 || bitslip_en_shift[1]==1'b0)begin
			bitslip_reg	<= 1'b0;
		end
		else begin
			if(bitslip_cnt==iv_line_length) begin	//ÿ�������ڼ��һ��ͬ����
				bitslip_reg	<= !data_lock;
			end
			else begin
				bitslip_reg	<= 1'b0;
			end
		end
	end
	assign	o_bitslip	= bitslip_reg	;

	//	===============================================================================================
	//	ref ***���***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	��������ź�
	//	-------------------------------------------------------------------------------------
	assign	o_data_valid	= data_lock;

	//	-------------------------------------------------------------------------------------
	//	������������ݣ����ִ�С��
	//	-------------------------------------------------------------------------------------
	genvar	l;
	generate
		for(l=0;l<CHANNEL_NUM;l=l+1) begin
			if(END_STYLE=="LITTLE") begin
				assign	ov_data[(l+1)*SENSOR_DAT_WIDTH-1:l*SENSOR_DAT_WIDTH]	= data_lane_align[l];
			end
			else if(END_STYLE=="BIG") begin
				assign	ov_data[(l+1)*SENSOR_DAT_WIDTH-1:l*SENSOR_DAT_WIDTH]	= data_lane_align[CHANNEL_NUM-l-1];
			end
		end
	endgenerate




endmodule