//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : harness
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/3/9 17:18:50	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------
`define		TESTCASE	testcase1
module harness ();

	//	ref signals
	//	===============================================================================================
	//	--ref parameter
	//	===============================================================================================
	parameter	FIFO_WIDTH	= `TESTCASE.FIFO_WIDTH	;
	parameter	FIFO_DEPTH	= `TESTCASE.FIFO_DEPTH	;

	//	===============================================================================================
	//	--ref signal
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	����
	//	-------------------------------------------------------------------------------------
	wire							reset_async	;
	wire							clk_wr	;
	wire							i_wr_en	;
	wire	[FIFO_WIDTH-1:0]		iv_fifo_din	;
	wire							clk_rd	;
	wire							i_rd_en	;

	//	-------------------------------------------------------------------------------------
	//	���
	//	-------------------------------------------------------------------------------------
	wire							o_fifo_full	;
	wire	[FIFO_WIDTH-1:0]		ov_fifo_dout	;
	wire							o_fifo_empty	;

	wire							full	;
	wire							empty	;
	wire	[7:0]					dout	;


	//	ref ARCHITECTURE

	//	-------------------------------------------------------------------------------------
	//	��������
	//	-------------------------------------------------------------------------------------
	assign	reset_async		= `TESTCASE.reset_async;
	assign	clk_wr			= `TESTCASE.clk_wr;
	assign	i_wr_en			= `TESTCASE.i_wr_en;
	assign	iv_fifo_din		= `TESTCASE.iv_fifo_din;
	assign	clk_rd			= `TESTCASE.clk_rd;
	assign	i_rd_en			= `TESTCASE.i_rd_en;

	//	-------------------------------------------------------------------------------------
	//	���� dut ģ��
	//	-------------------------------------------------------------------------------------
	async_fifo # (
	.FIFO_WIDTH		(FIFO_WIDTH		),
	.FIFO_DEPTH		(FIFO_DEPTH		)
	)
	async_fifo_inst (
	.reset_async	(reset_async	),
	.clk_wr			(clk_wr			),
	.i_wr_en		(i_wr_en		),
	.iv_fifo_din	(iv_fifo_din	),
	.o_fifo_full	(o_fifo_full	),
	.clk_rd			(clk_rd			),
	.i_rd_en		(i_rd_en		),
	.ov_fifo_dout	(ov_fifo_dout	),
	.o_fifo_empty	(o_fifo_empty	)
	);

	fifo_w8d16 fifo_w8d16_inst (
	.rst			(reset_async	),
	.wr_clk			(clk_wr			),
	.wr_en			(i_wr_en		),
	.full			(full			),
	.din			(iv_fifo_din	),
	.rd_clk			(clk_rd			),
	.rd_en			(i_rd_en		),
	.empty			(empty			),
	.dout			(dout			)
	);




	//generate vcd file
	//initial begin
	//$dumpfile("test.vcd");
	//$dumpvars(1,top_frame_buffer_inst);
	//end

	//for lattice simulation
	//GSR   GSR_INST (.GSR (1'b1)); //< global reset sig>
	//PUR   PUR_INST (.PUR (1'b1)); //<powerup reset sig>



endmodule
