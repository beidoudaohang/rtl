//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : counter
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2013/12/17 13:03:23	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------

//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

`timescale 1 ns / 1 ps
module counter (
	input 	 			clk		,		//ʱ��
	input				hend	,
	input 	 			i_clk_en,		//ʱ��ʹ��
	input 	 			i_aclr	,		//ͬ����λ
	output reg [15:0]	ov_q			//�������
	);

	always@(posedge clk) begin
		if(hend) begin
			if(i_aclr) begin
				ov_q <= 16'h0;
			end else if(i_clk_en) begin
				ov_q <= ov_q + 16'h1;
			end else begin
				ov_q <= ov_q;
			end
		end

	end

endmodule
