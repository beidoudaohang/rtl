//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : rd_back_buf
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/4/2 10:04:30	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module rd_back_buf # (
	parameter	DATA_WIDTH	= 8		//����λ��
	)
	(
	input						clk			,
	input						i_empty		,
	input	[DATA_WIDTH:0]		iv_pix_data	,
	output						o_rd		,
	output						o_fval		,
	output						o_lval		,
	output	[DATA_WIDTH-1:0]	ov_pix_data
	);

	//	ref signals


	//	ref ARCHITECTURE
	assign	o_rd		= !i_empty;
	assign	o_fval		= iv_pix_data[DATA_WIDTH];
	assign	o_lval		= o_fval&o_rd;
	assign	ov_pix_data	= iv_pix_data[DATA_WIDTH-1:0];
	


endmodule
