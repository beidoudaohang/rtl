//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : wb_gain
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/2/13 10:31:49	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ��ɫ��������ģ��
//              1)  : ������ʱ3��ʱ��
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module wb_gain # (
	parameter					SENSOR_DAT_WIDTH	= 10	,	//sensor ���ݿ��
	parameter					WB_GAIN_WIDTH		= 11	,	//��ƽ��ģ������Ĵ������
	parameter					WB_RATIO			= 8		,	//��ƽ��������ӣ��˷�������Ҫ���ƶ���λ
	parameter					REG_WD				= 32		//�Ĵ���λ��
	)
	(
	input								clk					,	//ʱ������
	input								i_fval				,	//���ź�
	input								i_lval				,	//���ź�
	input	[SENSOR_DAT_WIDTH-1:0]		iv_pix_data			,	//ͼ������
	input								i_r_flag			,	//��ɫ������־ R
	input								i_g_flag			,	//��ɫ������־ G
	input								i_b_flag			,	//��ɫ������־ B
	input	[REG_WD-1:0]				iv_pixel_format		,	//0x01080001:Mono8��0x01100003:Mono10��0x01080008:BayerGR8��0x0110000C:BayerGR10���ڰ׵�ʱ�򣬲����˷���
	input	[2:0]						iv_test_image_sel	,	//����ͼѡ��Ĵ���,000:��ʵͼ,001:����ͼ��1�Ҷ�ֵ֡����,110:����ͼ��2��ֹ��б����,010:����ͼ��3������б����
	input	[WB_GAIN_WIDTH-1:0]			iv_wb_gain_r		,	//��ƽ��R������R����С������256��Ľ����ȡֵ��Χ[0:2047]
	input	[WB_GAIN_WIDTH-1:0]			iv_wb_gain_g		,	//��ƽ��G������G����С������256��Ľ����ȡֵ��Χ[0:2047]
	input	[WB_GAIN_WIDTH-1:0]			iv_wb_gain_b		,	//��ƽ��B������B����С������256��Ľ����ȡֵ��Χ[0:2047]
	output								o_fval				,	//����Ч��o_fval��o_lval����λҪ��֤���������λһ��
	output								o_lval				,	//����Ч
	output	[SENSOR_DAT_WIDTH-1:0]		ov_pix_data				//ͼ������
	);

	//	ref signals
	reg														mono_sel		= 1'b0;
	wire													gain_enable		;
	reg		[WB_GAIN_WIDTH-1:0]								gain_coe		= {WB_GAIN_WIDTH{1'b0}};
	reg		[SENSOR_DAT_WIDTH-1:0]							pix_data_dly0	= {SENSOR_DAT_WIDTH{1'b0}};
	reg		[SENSOR_DAT_WIDTH-1:0]							pix_data_dly1	= {SENSOR_DAT_WIDTH{1'b0}};
	reg		[SENSOR_DAT_WIDTH-1:0]							pix_data_reg	= {SENSOR_DAT_WIDTH{1'b0}};
	wire	[16:0]											wb_mult_a		;
	wire	[16:0]											wb_mult_b		;
	wire	[33:0]											wb_mult_p		;
	reg														wb_mult_ce		= 1'b0;
	wire	[(WB_GAIN_WIDTH+SENSOR_DAT_WIDTH-1):0]			gain_all_data	;	//DSP�����������Ч������λ
	wire	[(WB_GAIN_WIDTH+SENSOR_DAT_WIDTH-WB_RATIO-1):0]	gain_reduce		;	//DSP�����������Ч������λ��λ֮��Ľ��
	wire	[(WB_GAIN_WIDTH-WB_RATIO-1):0]					gain_overflow	;	//DSP�����������Ч������λ�����λ
	reg														fval_dly0		= 1'b0;
	reg														fval_dly1		= 1'b0;
	reg														fval_dly2		= 1'b0;
	reg														lval_dly0		= 1'b0;
	reg														lval_dly1		= 1'b0;
	reg														lval_dly2		= 1'b0;
	reg		[WB_GAIN_WIDTH-1							:0]	wb_gain_r_m=0	;	//������Чʱ�����Ƶİ�ƽ����������
	reg		[WB_GAIN_WIDTH-1							:0]	wb_gain_g_m=0	;   //������Чʱ�����Ƶİ�ƽ������̷���
	reg		[WB_GAIN_WIDTH-1							:0]	wb_gain_b_m=0	;   //������Чʱ�����Ƶİ�ƽ�����������

	//	ref ARCHITECTURE
	//  ===============================================================================================
	//	ref ***��Чʱ��***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	���ظ�ʽѡ�кڰ�ģʽ
	//  -------------------------------------------------------------------------------------
	//  -------------------------------------------------------------------------------------
	//	Mono8		- 0x01080001	-> 0x1081	-> 0001,0000,1000,,,,0001
	//	Mono10		- 0x01100003	-> 0x1103	-> 0001,0001,0000,,,,0011
	//	BayerGR8	- 0x01080008	-> 0x1088	-> 0001,0000,1000,,,,1000
	//	BayerGR10	- 0x0110000C	-> 0x110C	-> 0001,0001,0000,,,,1100
	//											   --------!-!-------!!!!
	//                                                     ^    ^       ^------bit0
	//                                             bit20---|    |---bit16
	//	����� ! �ģ����ǲ���Ƚϵ�bit.�ֱ��� bit
	//  -------------------------------------------------------------------------------------
	//  -------------------------------------------------------------------------------------
	//	Ϊ�˱�����չ��ʹ��6bit�ж�����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		case({iv_pixel_format[20],iv_pixel_format[19],iv_pixel_format[3:0]})
			6'b010001	: mono_sel	<= 1'b1;
			6'b100011	: mono_sel	<= 1'b1;
			default		: mono_sel	<= 1'b0;
		endcase
	end

	//  -------------------------------------------------------------------------------------
	//	�˷�����ʹ�ܿ���
	//	1.�����ظ�ʽ�ǲ�ɫ����û��ѡ�в���ͼʱ���Ż����˷�����
	//	2.����ֱ���������
	//  -------------------------------------------------------------------------------------
	assign	gain_enable	= (mono_sel==1'b0 && iv_test_image_sel==3'b000) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//	����ϵ�� gain coefficient
	//  -------------------------------------------------------------------------------------

	always @ (posedge clk) begin
		if(!i_fval) begin
			wb_gain_r_m	<=  iv_wb_gain_r;
			wb_gain_g_m <=  iv_wb_gain_g;
			wb_gain_b_m <=  iv_wb_gain_b;
		end
	end

	always @ (posedge clk) begin
		if(i_r_flag) begin
			gain_coe	<= wb_gain_r_m;
		end
		else if(i_g_flag) begin
			gain_coe	<= wb_gain_g_m;
		end
		else if(i_b_flag) begin
			gain_coe	<= wb_gain_b_m;
		end
	end

	//  -------------------------------------------------------------------------------------
	//	������ʱ
	//	1.���� r g b �ı�־ѡ����ʵ����棬��Ҫ1��ʱ�䣬�������ҲҪ��ʱһ��
	//	2.DSP�˷�����ʱ1�ģ��������Ҫ��ʱ2�ģ�������DSP��������롣�Ա�����mux�߼���ѡ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		pix_data_dly0	<= iv_pix_data;
		pix_data_dly1	<= pix_data_dly0;
	end

	//  ===============================================================================================
	//	ref ***�˷������***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	�˷���
	//	1.ceʹ�ܣ�����������ݵ�ʱ��ʹ�ܹرգ���ʡ����
	//	2.�˷�������λ��17�����λ��34��Ŀ���Ƿ�����չ��DSP�ĸ�bitû���õ����ڲ��ֲ���ʱ�ᱻ�Ż���
	//	3.�ڲ���1��pipelin
	//  -------------------------------------------------------------------------------------
	wb_mult_a17b17p34 wb_mult_a17b17p34_inst (
	.clk	(clk		),
	.ce		(wb_mult_ce	),
	.a		(wb_mult_a	),
	.b		(wb_mult_b	),
	.p		(wb_mult_p	)
	);

	//  -------------------------------------------------------------------------------------
	//	�˷�����������˿�
	//	1.����˿ڶ���17bitλ��������������λ���㣬��Ҫ��0�����λ
	//	2.�˷���a��������ϵ��
	//	3.�˷���b������������
	//  -------------------------------------------------------------------------------------
	assign	wb_mult_a	= {{(17-WB_GAIN_WIDTH){1'b0}},gain_coe[WB_GAIN_WIDTH-1:0]};
	assign	wb_mult_b	= {{(17-SENSOR_DAT_WIDTH){1'b0}},pix_data_dly0[SENSOR_DAT_WIDTH-1:0]};

	//  -------------------------------------------------------------------------------------
	//	�˷���ʹ��
	//	1.������Чʹ��������ʹ�ܴ򿪵�ʱ�򣬳˷����Ż�ʹ��
	//	2.���򣬳˷���ʹ�ܹر�
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(gain_enable&i_lval) begin
			wb_mult_ce	<= 1'b1;
		end
		else begin
			wb_mult_ce	<= 1'b0;
		end
	end

	//  -------------------------------------------------------------------------------------
	//	���λ�Ľ���
	//	�˷�����������Ҫ���� WB_RATIO λ����Ϊ�˷�����ϵ����ʵ�ʵ�ϵ���ж�Ӧ��ϵ������ ����2λ���൱������ϵ����ʵ��ϵ����4����
	//  -------------------------------------------------------------------------------------
	//  -------------------------------------------------------------------------------------
	//	��������λ
	//	1.wb_mult_p		- �˷����ܹ�λ����34bit
	//	2.gain_all_data	- DSP��������ʵ����Чλ���� WB_GAIN_WIDTH + SENSOR_DAT_WIDTH����A�ڵĿ�� + B�ڵĿ�ȣ���λ��ȫ0
	//	3.gain_reduce	- DSP�������е���Ч����λ���� SENSOR_DAT_WIDTH + WB_RATIO�������а��������λ
	//	4.gain_overflow	- ���λ���� WB_GAIN_WIDTH + SENSOR_DAT_WIDTH - (SENSOR_DAT_WIDTH + WB_RATIO) = SENSOR_DAT_WIDTH - WB_RATIO
	//  -------------------------------------------------------------------------------------
	//	assign	gain_all_data	= wb_mult_p[(WB_GAIN_WIDTH+SENSOR_DAT_WIDTH-1):0];
	assign	gain_reduce		= wb_mult_p[(WB_GAIN_WIDTH+SENSOR_DAT_WIDTH-1):WB_RATIO];
	assign	gain_overflow	= wb_mult_p[(WB_GAIN_WIDTH+SENSOR_DAT_WIDTH-1):SENSOR_DAT_WIDTH+WB_RATIO];

	//  ===============================================================================================
	//	ref ***�������***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	�������������
	//	1.���г�����Чʱ
	//	--1.1���˷����治ʹ��ʱ��ֱ�������������ݡ�ʹ�ô�����֮������ݡ�
	//	--1.2���˷�����ʹ��ʱ��������λ��1���֣�˵���Ѿ����������Ч����Ϊȫ1
	//	--1.3���˷�����ʹ��ʱ�������λ��ȫ0���֣�˵��û�����������˷���������
	//	2.������ʱ����������Ϊ0
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(fval_dly1==1'b1 && lval_dly1==1'b1) begin
			if(!gain_enable) begin
				pix_data_reg	<= pix_data_dly1;
			end
			else begin
				if(|gain_overflow) begin
					pix_data_reg	<= {SENSOR_DAT_WIDTH{1'b1}};
				end
				else begin
					pix_data_reg	<= gain_reduce[SENSOR_DAT_WIDTH-1:0];
				end
			end
		end
		else begin
			pix_data_reg	<= {SENSOR_DAT_WIDTH{1'b0}};
		end
	end
	assign	ov_pix_data	= pix_data_reg;

	//  -------------------------------------------------------------------------------------
	//	�г��ź��ӳ� ���ӳ�3��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_dly0	<= i_fval;
		fval_dly1	<= fval_dly0;
		fval_dly2	<= fval_dly1;
	end
	assign	o_fval	= fval_dly2;

	//	-------------------------------------------------------------------------------------
	//	�����볡�ź�=0ʱ����������ź�Ҫ����
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		lval_dly0	<= i_lval;
		lval_dly1	<= lval_dly0;
		if(fval_dly1) begin
			lval_dly2	<= lval_dly1;
		end
		else begin
			lval_dly2	<= 1'b0;
		end
	end
	assign	o_lval	= lval_dly2;


endmodule