//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : bfm_sonyimx
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/4/3 15:04:32	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------
module bfm_sonyimx # (
	parameter	IMAGE_SRC				= "RANDOM"			,	//"RANDOM" or "FILE" or "LINE_INC" or "FRAME_INC" or "FRAME_INC_NO_RST"
	parameter	DATA_WIDTH				= 10				,	//���ݿ��
	parameter	SENSOR_CLK_DELAY_VALUE	= 0					,	//Sensor оƬ�ڲ���ʱ ��λns
	parameter	CLK_DATA_ALIGN			= "RISING"			,	//"RISING" - ���ʱ�ӵ������������ݶ��롣"FALLING" - ���ʱ�ӵ��½��������ݶ���
	parameter	FVAL_LVAL_ALIGN			= "FALSE"			,	//"TRUE" - fval �� lval ֮��ľ���̶�Ϊ3��ʱ�ӡ�"FALSE" - fval �� lval ֮��ľ��������趨
	parameter	SOURCE_FILE_PATH		= "source_file/"	,	//����Դ�ļ�·��
	parameter	GEN_FILE_EN				= 0					,	//0-���ɵ�ͼ��д���ļ���1-���ɵ�ͼ��д���ļ�
	parameter	GEN_FILE_PATH			= "gen_file/"		,	//����������Ҫд���·��
	parameter	NOISE_EN				= 0						//0-������������1-��������

	)
	(
	input		clk			,
	input		o_fval
	);

	//	ref signals
	//  -------------------------------------------------------------------------------------
	//	�������õļĴ���������
	//  -------------------------------------------------------------------------------------
	reg		[15:0]		iv_width					= 16'd16	;
	reg		[15:0]		iv_height					= 16'd16	;

	reg					reset		= 1'b0;
	reg					i_pause_en	= 1'b0;
	reg					i_continue_lval	= 1'b0;

	reg					pll_reset	= 1'b0;
	reg					data_init_done	= 1'b0;

	//	ref ARCHITECTURE

	//  ===============================================================================================
	//	ref ***task***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	--ref sensor pattern
	//  -------------------------------------------------------------------------------------
	task pattern_2para;
		input	[15:0]		width_input;
		input	[15:0]		height_input;
		begin
			#200
			iv_width			= width_input	;
			iv_height			= height_input	;
		end
	endtask


	//	-------------------------------------------------------------------------------------
	//	--ref sensor ��С��̬�л�
	//	-------------------------------------------------------------------------------------
	task pattern_random;
		input	[15:0]		start_point	;
		input	[15:0]		end_point	;

		reg		[15:0]		width;
		reg		[15:0]		height;
		begin
			//	-------------------------------------------------------------------------------------
			//	�� start point �� stop point ֮�䣬����һ�������.����8�ı���������2�ı�����
			//	-------------------------------------------------------------------------------------
			width	= $random()%(end_point-start_point)+start_point;
			width	= width+8-width%8;
			height	= $random()%(end_point-start_point)+start_point;
			height	= height+2-height%2;

			@ (negedge o_fval);
			reset	= 1'b1;
			@ (posedge clk);
			pattern_2para(width,height);
			@ (posedge clk);
			reset	= 1'b0;
		end
	endtask

	//	-------------------------------------------------------------------------------------
	//	--ref sensor ��λ
	//	-------------------------------------------------------------------------------------
	task reset_high;
		begin
			#1
			reset	= 1'b1;
		end
	endtask

	task reset_low;
		begin
			#1
			reset	= 1'b0;
		end
	endtask

	//	-------------------------------------------------------------------------------------
	//	ѭ����λsensor��ʹ֮������ͬ��С��ͼ��
	//	-------------------------------------------------------------------------------------
	task reset_repeat;
		integer		i;
		begin
			reset	= 1'b0;
			for(i=1;i<30;i=i+1) begin
				wait(o_fval==1'b1);
				repeat(i) @ (posedge clk);
				reset	= 1'b1;
				@ (posedge clk);
				reset	= 1'b0;
				repeat(20) @ (posedge clk);
			end
		end
	endtask

	//	-------------------------------------------------------------------------------------
	//	ѭ����λsensor��ʹ֮������ͬ��С��ͼ��
	//	-------------------------------------------------------------------------------------
	task reset_random;
		input	[15:0]		start_point	;
		input	[15:0]		end_point	;

		reg		[15:0]		time_slot;
		begin
			//	-------------------------------------------------------------------------------------
			//	�� start point �� stop point ֮�䣬����һ�������
			//	-------------------------------------------------------------------------------------
			time_slot	= $random()%(end_point-start_point)+start_point;
			@ (posedge o_fval);
			repeat(time_slot) @ (posedge clk);
			reset	= 1'b1;
			@ (posedge clk);
			reset	= 1'b0;
		end
	endtask

	//	-------------------------------------------------------------------------------------
	//	--ref pause_en ��ͣ
	//	-------------------------------------------------------------------------------------
	task pause_high;
		begin
			#1
			i_pause_en	= 1'b1;
		end
	endtask

	task pause_low;
		begin
			#1
			i_pause_en	= 1'b0;
		end
	endtask

	//	-------------------------------------------------------------------------------------
	//	--ref continue_lval ��ͣ
	//	-------------------------------------------------------------------------------------
	task continue_lval_high;
		begin
			#1
			i_continue_lval	= 1'b1;
		end
	endtask

	task continue_lval_low;
		begin
			#1
			i_continue_lval	= 1'b0;
		end
	endtask

	//	-------------------------------------------------------------------------------------
	//	--ref pll_reset
	//	-------------------------------------------------------------------------------------
	task pll_reset_high;
		begin
			#1
			pll_reset	= 1'b1;
		end
	endtask

	task pll_reset_low;
		begin
			#1
			pll_reset	= 1'b0;
		end
	endtask



endmodule
