//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : harness
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/3/9 17:18:50	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------
`define		TESTCASE	testcase_1
module harness ();

	//	ref signals
	//	===============================================================================================
	//	--ref parameter
	//	===============================================================================================
	parameter	FIFO_WIDTH	= `TESTCASE.FIFO_WIDTH		;
	parameter	FIFO_DEPTH	= `TESTCASE.FIFO_DEPTH		;

	//	===============================================================================================
	//	--ref signal
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	����
	//	-------------------------------------------------------------------------------------
	wire							reset		;
	wire							clk			;
	wire	[FIFO_WIDTH-1:0]		iv_din		;
	wire							i_wr		;
	wire							i_rd		;

	//	-------------------------------------------------------------------------------------
	//	���
	//	-------------------------------------------------------------------------------------
	wire							o_full		;
	wire							o_half_full	;
	wire							o_empty		;
	wire	[FIFO_WIDTH-1:0]		ov_dout		;

	//	-------------------------------------------------------------------------------------
	//	����
	//	-------------------------------------------------------------------------------------



	//	ref ARCHITECTURE

	//	-------------------------------------------------------------------------------------
	//	���������ź�
	//	-------------------------------------------------------------------------------------
	assign	clk						= `TESTCASE.clk		;
	assign	reset					= `TESTCASE.reset		;
	assign	iv_din					= `TESTCASE.iv_din	;
	assign	i_wr					= `TESTCASE.i_wr	;
	assign	i_rd					= `TESTCASE.i_rd	;


	//	-------------------------------------------------------------------------------------
	//	���� dut ģ��
	//	-------------------------------------------------------------------------------------
	sync_fifo_srl # (
	.FIFO_WIDTH		(FIFO_WIDTH	),
	.FIFO_DEPTH		(FIFO_DEPTH	)
	)
	sync_fifo_srl_inst (
	.reset			(reset			),
	.clk			(clk			),
	.iv_din			(iv_din			),
	.i_wr			(i_wr			),
	.o_full			(o_full			),
	.o_half_full	(o_half_full	),
	.i_rd			(i_rd			),
	.ov_dout		(ov_dout		),
	.o_empty		(o_empty		)
	);




	//generate vcd file
	//initial begin
	//$dumpfile("test.vcd");
	//$dumpvars(1,top_frame_buffer_inst);
	//end

	//for lattice simulation
	//GSR   GSR_INST (.GSR (1'b1)); //< global reset sig>
	//PUR   PUR_INST (.PUR (1'b1)); //<powerup reset sig>



endmodule
