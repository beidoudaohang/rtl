//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : wb_bayer_sel
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/2/13 10:22:58	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     : ����Sensor��bayer��ʽ����ֳ� R G B ������ɫ����
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module wb_bayer_sel # (
	parameter	BAYER_PATTERN		= "GR"	,	//"GR" "RG" "GB" "BG"
	parameter	SENSOR_DAT_WIDTH	= 10		//sensor ���ݿ��
	)
	(
	input								clk			,	//����ʱ��
	input								i_fval		,	//����Ч
	input								i_lval		,	//������Ч
	input	[SENSOR_DAT_WIDTH-1:0]		iv_pix_data	,	//ͼ������
	output								o_r_flag	,	//R ��־
	output								o_g_flag	,	//G ��־
	output								o_b_flag	,	//B ��־
	output								o_fval		,	//����Ч
	output								o_lval		,	//����Ч
	output	[SENSOR_DAT_WIDTH-1:0]		ov_pix_data		//ͼ������
	);

	//	ref signals
	reg									lval_dly		= 1'b0;
	wire								lval_fall		;
	reg									fval_dly		= 1'b0;
	reg		[SENSOR_DAT_WIDTH-1:0]		pix_data_dly	= {SENSOR_DAT_WIDTH{1'b0}};
	reg									line_cnt		= 1'b0;
	reg									r_flag			= 1'b0;
	reg									g_flag			= 1'b0;
	reg									b_flag			= 1'b0;

	//	ref ARCHITECTURE

	//  ===============================================================================================
	//	ref ***��ʱ ȡ����***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	����Чȡ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		lval_dly	<= i_lval;
	end
	assign	lval_fall	= (lval_dly==1'b1 && i_lval==1'b0) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//	��ʱ fval
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		fval_dly	<= i_fval;
	end

	//  -------------------------------------------------------------------------------------
	//	��ʱ pix data
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		pix_data_dly	<= iv_pix_data;
	end

	//  ===============================================================================================
	//	ref ***��ȡ��ɫ����***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	�м������������к�ż���е�bayer��ʽ��һ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!i_fval) begin
			line_cnt	<= 1'b0;
		end
		else begin
			if(lval_fall) begin
				line_cnt	<= !line_cnt;
			end
		end
	end

	//  -------------------------------------------------------------------------------------
	//	pattern �����ɫ����
	//  -------------------------------------------------------------------------------------
	generate
		//  -------------------------------------------------------------------------------------
		//	ref 1 GR pattern
		//	line 0		GRGRGRGR
		//		r flag	01010101
		//		g flag	10101010
		//		b flag	00000000
		//	line 1		BGBGBGBG
		//		r flag	00000000
		//		g flag	01010101
		//		b flag	10101010
		//  -------------------------------------------------------------------------------------
		if(BAYER_PATTERN=="GR") begin
			always @ (posedge clk) begin
				if(!i_lval) begin
					r_flag	<= 1'b0;
					g_flag	<= 1'b0;
					b_flag	<= 1'b0;
				end
				else begin
					if(!line_cnt) begin
						r_flag	<= g_flag;
						g_flag	<= !g_flag;
						b_flag	<= 1'b0;
					end
					else begin
						r_flag	<= 1'b0;
						g_flag	<= b_flag;
						b_flag	<= !b_flag;
					end
				end
			end
		end
		//  -------------------------------------------------------------------------------------
		//	ref 2 RG pattern
		//	line 0		RGRGRGRG
		//		r flag	10101010
		//		g flag	01010101
		//		b flag	00000000
		//	line 1		GBGBGBGB
		//		r flag	00000000
		//		g flag	10101010
		//		b flag	01010101
		//  -------------------------------------------------------------------------------------
		else if(BAYER_PATTERN=="RG") begin
			always @ (posedge clk) begin
				if(!i_lval) begin
					r_flag	<= 1'b0;
					g_flag	<= 1'b0;
					b_flag	<= 1'b0;
				end
				else begin
					if(!line_cnt) begin
						r_flag	<= !r_flag;
						g_flag	<= r_flag;
						b_flag	<= 1'b0;
					end
					else begin
						r_flag	<= 1'b0;
						g_flag	<= !g_flag;
						b_flag	<= g_flag;
					end
				end
			end
		end
		//  -------------------------------------------------------------------------------------
		//	ref 3 GB pattern
		//	line 0		GBGBGBGB
		//		r flag	00000000
		//		g flag	10101010
		//		b flag	01010101
		//	line 1		RGRGRGRG
		//		r flag	10101010
		//		g flag	01010101
		//		b flag	00000000
		//  -------------------------------------------------------------------------------------
		else if(BAYER_PATTERN=="GB") begin
			always @ (posedge clk) begin
				if(!i_lval) begin
					r_flag	<= 1'b0;
					g_flag	<= 1'b0;
					b_flag	<= 1'b0;
				end
				else begin
					if(!line_cnt) begin
						r_flag	<= 1'b0;
						g_flag	<= !g_flag;
						b_flag	<= g_flag;
					end
					else begin
						r_flag	<= !r_flag;
						g_flag	<= r_flag;
						b_flag	<= 1'b0;
					end
				end
			end
		end
		//  -------------------------------------------------------------------------------------
		//	ref 4 BG pattern
		//	line 0		BGBGBGBG
		//		r flag	00000000
		//		g flag	01010101
		//		b flag	10101010
		//	line 1		GRGRGRGR
		//		r flag	01010101
		//		g flag	10101010
		//		b flag	00000000
		//  -------------------------------------------------------------------------------------
		else if(BAYER_PATTERN=="BG") begin
			always @ (posedge clk) begin
				if(!i_lval) begin
					r_flag	<= 1'b0;
					g_flag	<= 1'b0;
					b_flag	<= 1'b0;
				end
				else begin
					if(!line_cnt) begin
						r_flag	<= 1'b0;
						g_flag	<= b_flag;
						b_flag	<= !b_flag;
					end
					else begin
						r_flag	<= g_flag;
						g_flag	<= !g_flag;
						b_flag	<= 1'b0;
					end
				end
			end
		end
		//  -------------------------------------------------------------------------------------
		//	���������Ĳ���������
		//  -------------------------------------------------------------------------------------
		else begin
			always @ (posedge clk) begin
				r_flag	<= 1'b0;
				g_flag	<= 1'b0;
				b_flag	<= 1'b0;
			end
		end

	endgenerate

	//  -------------------------------------------------------------------------------------
	//	�����ɫ������־
	//  -------------------------------------------------------------------------------------
	assign	o_r_flag	= r_flag;
	assign	o_g_flag	= g_flag;
	assign	o_b_flag	= b_flag;

	//  ===============================================================================================
	//	ref ***�����������***
	//  ===============================================================================================
	assign	o_fval		= 	fval_dly;
	assign	o_lval		= 	lval_dly;
	assign	ov_pix_data	= 	pix_data_dly;










endmodule
